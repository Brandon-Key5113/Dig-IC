
--
-- Definition of  Multiplier
--
--      Sun Nov 17 16:34:50 2019
--
--      LeonardoSpectrum Level 3, 2008b.3
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library gdk;
use gdk.gdk_comps.all;

entity Multiplier is
   port (
      A : IN std_logic_vector (15 DOWNTO 0) ;
      B : IN std_logic_vector (15 DOWNTO 0) ;
      Product : OUT std_logic_vector (31 DOWNTO 0)) ;
end Multiplier ;

architecture Behavioral of Multiplier is
   component FA_1bit
      port (
         A : IN std_logic ;
         B : IN std_logic ;
         Cin : IN std_logic ;
         S : OUT std_logic ;
         Cout : OUT std_logic) ;
   end component ;
   signal F_239, F_238, F_237, F_236, F_235, F_234, F_233, F_232, F_231,
      F_230, F_229, F_228, F_227, F_226, F_225, F_223, F_222, F_221, F_220,
      F_219, F_218, F_217, F_216, F_215, F_214, F_213, F_212, F_211, F_210,
      F_209, F_207, F_206, F_205, F_204, F_203, F_202, F_201, F_200, F_199,
      F_198, F_197, F_196, F_195, F_194, F_193, F_191, F_190, F_189, F_188,
      F_187, F_186, F_185, F_184, F_183, F_182, F_181, F_180, F_179, F_178,
      F_177, F_175, F_174, F_173, F_172, F_171, F_170, F_169, F_168, F_167,
      F_166, F_165, F_164, F_163, F_162, F_161, F_159, F_158, F_157, F_156,
      F_155, F_154, F_153, F_152, F_151, F_150, F_149, F_148, F_147, F_146,
      F_145, F_143, F_142, F_141, F_140, F_139, F_138, F_137, F_136, F_135,
      F_134, F_133, F_132, F_131, F_130, F_129, F_127, F_126, F_125, F_124,
      F_123, F_122, F_121, F_120, F_119, F_118, F_117, F_116, F_115, F_114,
      F_113, F_111, F_110, F_109, F_108, F_107, F_106, F_105, F_104, F_103,
      F_102, F_101, F_100, F_99, F_98, F_97, F_95, F_94, F_93, F_92, F_91,
      F_90, F_89, F_88, F_87, F_86, F_85, F_84, F_83, F_82, F_81, F_79, F_78,
      F_77, F_76, F_75, F_74, F_73, F_72, F_71, F_70, F_69, F_68, F_67, F_66,
      F_65, F_63, F_62, F_61, F_60, F_59, F_58, F_57, F_56, F_55, F_54, F_53,
      F_52, F_51, F_50, F_49, F_47, F_46, F_45, F_44, F_43, F_42, F_41, F_40,
      F_39, F_38, F_37, F_36, F_35, F_34, F_33, F_31, F_30, F_29, F_28, F_27,
      F_26, F_25, F_24, F_23, F_22, F_21, F_20, F_19, F_18, F_17, F_15, F_14,
      F_13, F_12, F_11, F_10, F_9, F_8, F_7, F_6, F_5, F_4, F_3, F_2, F_1,
      CoutArray_254, CoutArray_253, CoutArray_252, CoutArray_251,
      CoutArray_250, CoutArray_249, CoutArray_248, CoutArray_247,
      CoutArray_246, CoutArray_245, CoutArray_244, CoutArray_243,
      CoutArray_242, CoutArray_241, CoutArray_240, CoutArray_239,
      CoutArray_238, CoutArray_237, CoutArray_236, CoutArray_235,
      CoutArray_234, CoutArray_233, CoutArray_232, CoutArray_231,
      CoutArray_230, CoutArray_229, CoutArray_228, CoutArray_227,
      CoutArray_226, CoutArray_225, CoutArray_224, CoutArray_223,
      CoutArray_222, CoutArray_221, CoutArray_220, CoutArray_219,
      CoutArray_218, CoutArray_217, CoutArray_216, CoutArray_215,
      CoutArray_214, CoutArray_213, CoutArray_212, CoutArray_211,
      CoutArray_210, CoutArray_209, CoutArray_208, CoutArray_207,
      CoutArray_206, CoutArray_205, CoutArray_204, CoutArray_203,
      CoutArray_202, CoutArray_201, CoutArray_200, CoutArray_199,
      CoutArray_198, CoutArray_197, CoutArray_196, CoutArray_195,
      CoutArray_194, CoutArray_193, CoutArray_192, CoutArray_191,
      CoutArray_190, CoutArray_189, CoutArray_188, CoutArray_187,
      CoutArray_186, CoutArray_185, CoutArray_184, CoutArray_183,
      CoutArray_182, CoutArray_181, CoutArray_180, CoutArray_179,
      CoutArray_178, CoutArray_177, CoutArray_176, CoutArray_175,
      CoutArray_174, CoutArray_173, CoutArray_172, CoutArray_171,
      CoutArray_170, CoutArray_169, CoutArray_168, CoutArray_167,
      CoutArray_166, CoutArray_165, CoutArray_164, CoutArray_163,
      CoutArray_162, CoutArray_161, CoutArray_160, CoutArray_159,
      CoutArray_158, CoutArray_157, CoutArray_156, CoutArray_155,
      CoutArray_154, CoutArray_153, CoutArray_152, CoutArray_151,
      CoutArray_150, CoutArray_149, CoutArray_148, CoutArray_147,
      CoutArray_146, CoutArray_145, CoutArray_144, CoutArray_143,
      CoutArray_142, CoutArray_141, CoutArray_140, CoutArray_139,
      CoutArray_138, CoutArray_137, CoutArray_136, CoutArray_135,
      CoutArray_134, CoutArray_133, CoutArray_132, CoutArray_131,
      CoutArray_130, CoutArray_129, CoutArray_128, CoutArray_127,
      CoutArray_126, CoutArray_125, CoutArray_124, CoutArray_123,
      CoutArray_122, CoutArray_121, CoutArray_120, CoutArray_119,
      CoutArray_118, CoutArray_117, CoutArray_116, CoutArray_115,
      CoutArray_114, CoutArray_113, CoutArray_112, CoutArray_111,
      CoutArray_110, CoutArray_109, CoutArray_108, CoutArray_107,
      CoutArray_106, CoutArray_105, CoutArray_104, CoutArray_103,
      CoutArray_102, CoutArray_101, CoutArray_100, CoutArray_99,
      CoutArray_98, CoutArray_97, CoutArray_96, CoutArray_95, CoutArray_94,
      CoutArray_93, CoutArray_92, CoutArray_91, CoutArray_90, CoutArray_89,
      CoutArray_88, CoutArray_87, CoutArray_86, CoutArray_85, CoutArray_84,
      CoutArray_83, CoutArray_82, CoutArray_81, CoutArray_80, CoutArray_79,
      CoutArray_78, CoutArray_77, CoutArray_76, CoutArray_75, CoutArray_74,
      CoutArray_73, CoutArray_72, CoutArray_71, CoutArray_70, CoutArray_69,
      CoutArray_68, CoutArray_67, CoutArray_66, CoutArray_65, CoutArray_64,
      CoutArray_63, CoutArray_62, CoutArray_61, CoutArray_60, CoutArray_59,
      CoutArray_58, CoutArray_57, CoutArray_56, CoutArray_55, CoutArray_54,
      CoutArray_53, CoutArray_52, CoutArray_51, CoutArray_50, CoutArray_49,
      CoutArray_48, CoutArray_47, CoutArray_46, CoutArray_45, CoutArray_44,
      CoutArray_43, CoutArray_42, CoutArray_41, CoutArray_40, CoutArray_39,
      CoutArray_38, CoutArray_37, CoutArray_36, CoutArray_35, CoutArray_34,
      CoutArray_33, CoutArray_32, CoutArray_31, CoutArray_30, CoutArray_29,
      CoutArray_28, CoutArray_27, CoutArray_26, CoutArray_25, CoutArray_24,
      CoutArray_23, CoutArray_22, CoutArray_21, CoutArray_20, CoutArray_19,
      CoutArray_18, CoutArray_17, CoutArray_16,
      forrow_1_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_1_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_1_ifn0_forcol_15_GEN1N_ANDADD1N_F,
      forrow_2_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_2_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_2_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_3_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_3_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_3_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_4_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_4_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_4_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_5_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_5_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_5_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_6_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_6_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_6_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_7_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_7_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_7_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_8_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_8_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_8_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_9_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_9_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_9_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_10_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_10_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_10_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_11_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_11_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_11_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_12_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_12_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_12_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_13_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_13_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_13_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_14_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_14_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_14_ifn0_forcol_15_GENN_ANDADDN_F,
      forrow_15_ifn0_forcol_0_GEN0_ANDADD0_F,
      forrow_15_ifn0_forcol_1_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_2_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_3_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_4_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_5_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_6_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_7_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_8_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_9_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_10_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_11_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_12_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_13_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_14_GENX_ANDADDX_F,
      forrow_15_ifn0_forcol_15_GENN_ANDADDN_F, F_1024: std_logic ;

begin
   forrow_1_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_1, Cin=>F_1024, S=>
      Product(1), Cout=>CoutArray_16);
   forrow_1_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_2, Cin=>CoutArray_16, S=>
      F_17, Cout=>CoutArray_17);
   forrow_1_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_3, Cin=>CoutArray_17, S=>
      F_18, Cout=>CoutArray_18);
   forrow_1_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_4, Cin=>CoutArray_18, S=>
      F_19, Cout=>CoutArray_19);
   forrow_1_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_5, Cin=>CoutArray_19, S=>
      F_20, Cout=>CoutArray_20);
   forrow_1_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_6, Cin=>CoutArray_20, S=>
      F_21, Cout=>CoutArray_21);
   forrow_1_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_7, Cin=>CoutArray_21, S=>
      F_22, Cout=>CoutArray_22);
   forrow_1_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_8, Cin=>CoutArray_22, S=>
      F_23, Cout=>CoutArray_23);
   forrow_1_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_9, Cin=>CoutArray_23, S=>
      F_24, Cout=>CoutArray_24);
   forrow_1_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_10, Cin=>CoutArray_24, S=>
      F_25, Cout=>CoutArray_25);
   forrow_1_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_11, Cin=>CoutArray_25, S
      =>F_26, Cout=>CoutArray_26);
   forrow_1_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_12, Cin=>CoutArray_26, S
      =>F_27, Cout=>CoutArray_27);
   forrow_1_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_13, Cin=>CoutArray_27, S
      =>F_28, Cout=>CoutArray_28);
   forrow_1_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_14, Cin=>CoutArray_28, S
      =>F_29, Cout=>CoutArray_29);
   forrow_1_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_15, Cin=>CoutArray_29, S
      =>F_30, Cout=>CoutArray_30);
   forrow_1_ifn0_forcol_15_GEN1N_ANDADD1N_FA : FA_1bit port map ( A=>
      forrow_1_ifn0_forcol_15_GEN1N_ANDADD1N_F, B=>F_1024, Cin=>CoutArray_30,
      S=>F_31, Cout=>CoutArray_31);
   forrow_2_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_17, Cin=>F_1024, S=>
      Product(2), Cout=>CoutArray_32);
   forrow_2_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_18, Cin=>CoutArray_32, S=>
      F_33, Cout=>CoutArray_33);
   forrow_2_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_19, Cin=>CoutArray_33, S=>
      F_34, Cout=>CoutArray_34);
   forrow_2_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_20, Cin=>CoutArray_34, S=>
      F_35, Cout=>CoutArray_35);
   forrow_2_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_21, Cin=>CoutArray_35, S=>
      F_36, Cout=>CoutArray_36);
   forrow_2_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_22, Cin=>CoutArray_36, S=>
      F_37, Cout=>CoutArray_37);
   forrow_2_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_23, Cin=>CoutArray_37, S=>
      F_38, Cout=>CoutArray_38);
   forrow_2_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_24, Cin=>CoutArray_38, S=>
      F_39, Cout=>CoutArray_39);
   forrow_2_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_25, Cin=>CoutArray_39, S=>
      F_40, Cout=>CoutArray_40);
   forrow_2_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_26, Cin=>CoutArray_40, S=>
      F_41, Cout=>CoutArray_41);
   forrow_2_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_27, Cin=>CoutArray_41, S
      =>F_42, Cout=>CoutArray_42);
   forrow_2_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_28, Cin=>CoutArray_42, S
      =>F_43, Cout=>CoutArray_43);
   forrow_2_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_29, Cin=>CoutArray_43, S
      =>F_44, Cout=>CoutArray_44);
   forrow_2_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_30, Cin=>CoutArray_44, S
      =>F_45, Cout=>CoutArray_45);
   forrow_2_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_31, Cin=>CoutArray_45, S
      =>F_46, Cout=>CoutArray_46);
   forrow_2_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_2_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_31, Cin=>
      CoutArray_46, S=>F_47, Cout=>CoutArray_47);
   forrow_3_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_33, Cin=>F_1024, S=>
      Product(3), Cout=>CoutArray_48);
   forrow_3_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_34, Cin=>CoutArray_48, S=>
      F_49, Cout=>CoutArray_49);
   forrow_3_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_35, Cin=>CoutArray_49, S=>
      F_50, Cout=>CoutArray_50);
   forrow_3_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_36, Cin=>CoutArray_50, S=>
      F_51, Cout=>CoutArray_51);
   forrow_3_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_37, Cin=>CoutArray_51, S=>
      F_52, Cout=>CoutArray_52);
   forrow_3_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_38, Cin=>CoutArray_52, S=>
      F_53, Cout=>CoutArray_53);
   forrow_3_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_39, Cin=>CoutArray_53, S=>
      F_54, Cout=>CoutArray_54);
   forrow_3_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_40, Cin=>CoutArray_54, S=>
      F_55, Cout=>CoutArray_55);
   forrow_3_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_41, Cin=>CoutArray_55, S=>
      F_56, Cout=>CoutArray_56);
   forrow_3_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_42, Cin=>CoutArray_56, S=>
      F_57, Cout=>CoutArray_57);
   forrow_3_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_43, Cin=>CoutArray_57, S
      =>F_58, Cout=>CoutArray_58);
   forrow_3_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_44, Cin=>CoutArray_58, S
      =>F_59, Cout=>CoutArray_59);
   forrow_3_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_45, Cin=>CoutArray_59, S
      =>F_60, Cout=>CoutArray_60);
   forrow_3_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_46, Cin=>CoutArray_60, S
      =>F_61, Cout=>CoutArray_61);
   forrow_3_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_47, Cin=>CoutArray_61, S
      =>F_62, Cout=>CoutArray_62);
   forrow_3_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_3_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_47, Cin=>
      CoutArray_62, S=>F_63, Cout=>CoutArray_63);
   forrow_4_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_49, Cin=>F_1024, S=>
      Product(4), Cout=>CoutArray_64);
   forrow_4_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_50, Cin=>CoutArray_64, S=>
      F_65, Cout=>CoutArray_65);
   forrow_4_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_51, Cin=>CoutArray_65, S=>
      F_66, Cout=>CoutArray_66);
   forrow_4_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_52, Cin=>CoutArray_66, S=>
      F_67, Cout=>CoutArray_67);
   forrow_4_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_53, Cin=>CoutArray_67, S=>
      F_68, Cout=>CoutArray_68);
   forrow_4_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_54, Cin=>CoutArray_68, S=>
      F_69, Cout=>CoutArray_69);
   forrow_4_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_55, Cin=>CoutArray_69, S=>
      F_70, Cout=>CoutArray_70);
   forrow_4_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_56, Cin=>CoutArray_70, S=>
      F_71, Cout=>CoutArray_71);
   forrow_4_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_57, Cin=>CoutArray_71, S=>
      F_72, Cout=>CoutArray_72);
   forrow_4_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_58, Cin=>CoutArray_72, S=>
      F_73, Cout=>CoutArray_73);
   forrow_4_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_59, Cin=>CoutArray_73, S
      =>F_74, Cout=>CoutArray_74);
   forrow_4_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_60, Cin=>CoutArray_74, S
      =>F_75, Cout=>CoutArray_75);
   forrow_4_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_61, Cin=>CoutArray_75, S
      =>F_76, Cout=>CoutArray_76);
   forrow_4_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_62, Cin=>CoutArray_76, S
      =>F_77, Cout=>CoutArray_77);
   forrow_4_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_63, Cin=>CoutArray_77, S
      =>F_78, Cout=>CoutArray_78);
   forrow_4_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_4_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_63, Cin=>
      CoutArray_78, S=>F_79, Cout=>CoutArray_79);
   forrow_5_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_65, Cin=>F_1024, S=>
      Product(5), Cout=>CoutArray_80);
   forrow_5_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_66, Cin=>CoutArray_80, S=>
      F_81, Cout=>CoutArray_81);
   forrow_5_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_67, Cin=>CoutArray_81, S=>
      F_82, Cout=>CoutArray_82);
   forrow_5_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_68, Cin=>CoutArray_82, S=>
      F_83, Cout=>CoutArray_83);
   forrow_5_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_69, Cin=>CoutArray_83, S=>
      F_84, Cout=>CoutArray_84);
   forrow_5_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_70, Cin=>CoutArray_84, S=>
      F_85, Cout=>CoutArray_85);
   forrow_5_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_71, Cin=>CoutArray_85, S=>
      F_86, Cout=>CoutArray_86);
   forrow_5_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_72, Cin=>CoutArray_86, S=>
      F_87, Cout=>CoutArray_87);
   forrow_5_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_73, Cin=>CoutArray_87, S=>
      F_88, Cout=>CoutArray_88);
   forrow_5_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_74, Cin=>CoutArray_88, S=>
      F_89, Cout=>CoutArray_89);
   forrow_5_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_75, Cin=>CoutArray_89, S
      =>F_90, Cout=>CoutArray_90);
   forrow_5_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_76, Cin=>CoutArray_90, S
      =>F_91, Cout=>CoutArray_91);
   forrow_5_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_77, Cin=>CoutArray_91, S
      =>F_92, Cout=>CoutArray_92);
   forrow_5_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_78, Cin=>CoutArray_92, S
      =>F_93, Cout=>CoutArray_93);
   forrow_5_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_79, Cin=>CoutArray_93, S
      =>F_94, Cout=>CoutArray_94);
   forrow_5_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_5_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_79, Cin=>
      CoutArray_94, S=>F_95, Cout=>CoutArray_95);
   forrow_6_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_81, Cin=>F_1024, S=>
      Product(6), Cout=>CoutArray_96);
   forrow_6_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_82, Cin=>CoutArray_96, S=>
      F_97, Cout=>CoutArray_97);
   forrow_6_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_83, Cin=>CoutArray_97, S=>
      F_98, Cout=>CoutArray_98);
   forrow_6_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_84, Cin=>CoutArray_98, S=>
      F_99, Cout=>CoutArray_99);
   forrow_6_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_85, Cin=>CoutArray_99, S=>
      F_100, Cout=>CoutArray_100);
   forrow_6_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_86, Cin=>CoutArray_100, S
      =>F_101, Cout=>CoutArray_101);
   forrow_6_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_87, Cin=>CoutArray_101, S
      =>F_102, Cout=>CoutArray_102);
   forrow_6_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_88, Cin=>CoutArray_102, S
      =>F_103, Cout=>CoutArray_103);
   forrow_6_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_89, Cin=>CoutArray_103, S
      =>F_104, Cout=>CoutArray_104);
   forrow_6_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_90, Cin=>CoutArray_104, S
      =>F_105, Cout=>CoutArray_105);
   forrow_6_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_91, Cin=>CoutArray_105, S
      =>F_106, Cout=>CoutArray_106);
   forrow_6_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_92, Cin=>CoutArray_106, S
      =>F_107, Cout=>CoutArray_107);
   forrow_6_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_93, Cin=>CoutArray_107, S
      =>F_108, Cout=>CoutArray_108);
   forrow_6_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_94, Cin=>CoutArray_108, S
      =>F_109, Cout=>CoutArray_109);
   forrow_6_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_95, Cin=>CoutArray_109, S
      =>F_110, Cout=>CoutArray_110);
   forrow_6_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_6_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_95, Cin=>
      CoutArray_110, S=>F_111, Cout=>CoutArray_111);
   forrow_7_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_97, Cin=>F_1024, S=>
      Product(7), Cout=>CoutArray_112);
   forrow_7_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_98, Cin=>CoutArray_112, S
      =>F_113, Cout=>CoutArray_113);
   forrow_7_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_99, Cin=>CoutArray_113, S
      =>F_114, Cout=>CoutArray_114);
   forrow_7_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_100, Cin=>CoutArray_114, S
      =>F_115, Cout=>CoutArray_115);
   forrow_7_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_101, Cin=>CoutArray_115, S
      =>F_116, Cout=>CoutArray_116);
   forrow_7_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_102, Cin=>CoutArray_116, S
      =>F_117, Cout=>CoutArray_117);
   forrow_7_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_103, Cin=>CoutArray_117, S
      =>F_118, Cout=>CoutArray_118);
   forrow_7_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_104, Cin=>CoutArray_118, S
      =>F_119, Cout=>CoutArray_119);
   forrow_7_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_105, Cin=>CoutArray_119, S
      =>F_120, Cout=>CoutArray_120);
   forrow_7_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_106, Cin=>CoutArray_120, S
      =>F_121, Cout=>CoutArray_121);
   forrow_7_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_107, Cin=>CoutArray_121,
      S=>F_122, Cout=>CoutArray_122);
   forrow_7_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_108, Cin=>CoutArray_122,
      S=>F_123, Cout=>CoutArray_123);
   forrow_7_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_109, Cin=>CoutArray_123,
      S=>F_124, Cout=>CoutArray_124);
   forrow_7_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_110, Cin=>CoutArray_124,
      S=>F_125, Cout=>CoutArray_125);
   forrow_7_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_111, Cin=>CoutArray_125,
      S=>F_126, Cout=>CoutArray_126);
   forrow_7_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_7_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_111, Cin=>
      CoutArray_126, S=>F_127, Cout=>CoutArray_127);
   forrow_8_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_113, Cin=>F_1024, S=>
      Product(8), Cout=>CoutArray_128);
   forrow_8_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_114, Cin=>CoutArray_128, S
      =>F_129, Cout=>CoutArray_129);
   forrow_8_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_115, Cin=>CoutArray_129, S
      =>F_130, Cout=>CoutArray_130);
   forrow_8_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_116, Cin=>CoutArray_130, S
      =>F_131, Cout=>CoutArray_131);
   forrow_8_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_117, Cin=>CoutArray_131, S
      =>F_132, Cout=>CoutArray_132);
   forrow_8_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_118, Cin=>CoutArray_132, S
      =>F_133, Cout=>CoutArray_133);
   forrow_8_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_119, Cin=>CoutArray_133, S
      =>F_134, Cout=>CoutArray_134);
   forrow_8_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_120, Cin=>CoutArray_134, S
      =>F_135, Cout=>CoutArray_135);
   forrow_8_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_121, Cin=>CoutArray_135, S
      =>F_136, Cout=>CoutArray_136);
   forrow_8_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_122, Cin=>CoutArray_136, S
      =>F_137, Cout=>CoutArray_137);
   forrow_8_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_123, Cin=>CoutArray_137,
      S=>F_138, Cout=>CoutArray_138);
   forrow_8_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_124, Cin=>CoutArray_138,
      S=>F_139, Cout=>CoutArray_139);
   forrow_8_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_125, Cin=>CoutArray_139,
      S=>F_140, Cout=>CoutArray_140);
   forrow_8_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_126, Cin=>CoutArray_140,
      S=>F_141, Cout=>CoutArray_141);
   forrow_8_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_127, Cin=>CoutArray_141,
      S=>F_142, Cout=>CoutArray_142);
   forrow_8_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_8_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_127, Cin=>
      CoutArray_142, S=>F_143, Cout=>CoutArray_143);
   forrow_9_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_129, Cin=>F_1024, S=>
      Product(9), Cout=>CoutArray_144);
   forrow_9_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_130, Cin=>CoutArray_144, S
      =>F_145, Cout=>CoutArray_145);
   forrow_9_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_131, Cin=>CoutArray_145, S
      =>F_146, Cout=>CoutArray_146);
   forrow_9_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_132, Cin=>CoutArray_146, S
      =>F_147, Cout=>CoutArray_147);
   forrow_9_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_133, Cin=>CoutArray_147, S
      =>F_148, Cout=>CoutArray_148);
   forrow_9_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_134, Cin=>CoutArray_148, S
      =>F_149, Cout=>CoutArray_149);
   forrow_9_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_135, Cin=>CoutArray_149, S
      =>F_150, Cout=>CoutArray_150);
   forrow_9_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_136, Cin=>CoutArray_150, S
      =>F_151, Cout=>CoutArray_151);
   forrow_9_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_137, Cin=>CoutArray_151, S
      =>F_152, Cout=>CoutArray_152);
   forrow_9_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_138, Cin=>CoutArray_152, S
      =>F_153, Cout=>CoutArray_153);
   forrow_9_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_139, Cin=>CoutArray_153,
      S=>F_154, Cout=>CoutArray_154);
   forrow_9_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_140, Cin=>CoutArray_154,
      S=>F_155, Cout=>CoutArray_155);
   forrow_9_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_141, Cin=>CoutArray_155,
      S=>F_156, Cout=>CoutArray_156);
   forrow_9_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_142, Cin=>CoutArray_156,
      S=>F_157, Cout=>CoutArray_157);
   forrow_9_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_143, Cin=>CoutArray_157,
      S=>F_158, Cout=>CoutArray_158);
   forrow_9_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_9_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_143, Cin=>
      CoutArray_158, S=>F_159, Cout=>CoutArray_159);
   forrow_10_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_145, Cin=>F_1024, S=>
      Product(10), Cout=>CoutArray_160);
   forrow_10_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_146, Cin=>CoutArray_160,
      S=>F_161, Cout=>CoutArray_161);
   forrow_10_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_147, Cin=>CoutArray_161,
      S=>F_162, Cout=>CoutArray_162);
   forrow_10_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_148, Cin=>CoutArray_162,
      S=>F_163, Cout=>CoutArray_163);
   forrow_10_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_149, Cin=>CoutArray_163,
      S=>F_164, Cout=>CoutArray_164);
   forrow_10_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_150, Cin=>CoutArray_164,
      S=>F_165, Cout=>CoutArray_165);
   forrow_10_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_151, Cin=>CoutArray_165,
      S=>F_166, Cout=>CoutArray_166);
   forrow_10_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_152, Cin=>CoutArray_166,
      S=>F_167, Cout=>CoutArray_167);
   forrow_10_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_153, Cin=>CoutArray_167,
      S=>F_168, Cout=>CoutArray_168);
   forrow_10_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_154, Cin=>CoutArray_168,
      S=>F_169, Cout=>CoutArray_169);
   forrow_10_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_155, Cin=>CoutArray_169,
      S=>F_170, Cout=>CoutArray_170);
   forrow_10_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_156, Cin=>CoutArray_170,
      S=>F_171, Cout=>CoutArray_171);
   forrow_10_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_157, Cin=>CoutArray_171,
      S=>F_172, Cout=>CoutArray_172);
   forrow_10_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_158, Cin=>CoutArray_172,
      S=>F_173, Cout=>CoutArray_173);
   forrow_10_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_159, Cin=>CoutArray_173,
      S=>F_174, Cout=>CoutArray_174);
   forrow_10_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_10_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_159, Cin=>
      CoutArray_174, S=>F_175, Cout=>CoutArray_175);
   forrow_11_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_161, Cin=>F_1024, S=>
      Product(11), Cout=>CoutArray_176);
   forrow_11_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_162, Cin=>CoutArray_176,
      S=>F_177, Cout=>CoutArray_177);
   forrow_11_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_163, Cin=>CoutArray_177,
      S=>F_178, Cout=>CoutArray_178);
   forrow_11_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_164, Cin=>CoutArray_178,
      S=>F_179, Cout=>CoutArray_179);
   forrow_11_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_165, Cin=>CoutArray_179,
      S=>F_180, Cout=>CoutArray_180);
   forrow_11_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_166, Cin=>CoutArray_180,
      S=>F_181, Cout=>CoutArray_181);
   forrow_11_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_167, Cin=>CoutArray_181,
      S=>F_182, Cout=>CoutArray_182);
   forrow_11_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_168, Cin=>CoutArray_182,
      S=>F_183, Cout=>CoutArray_183);
   forrow_11_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_169, Cin=>CoutArray_183,
      S=>F_184, Cout=>CoutArray_184);
   forrow_11_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_170, Cin=>CoutArray_184,
      S=>F_185, Cout=>CoutArray_185);
   forrow_11_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_171, Cin=>CoutArray_185,
      S=>F_186, Cout=>CoutArray_186);
   forrow_11_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_172, Cin=>CoutArray_186,
      S=>F_187, Cout=>CoutArray_187);
   forrow_11_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_173, Cin=>CoutArray_187,
      S=>F_188, Cout=>CoutArray_188);
   forrow_11_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_174, Cin=>CoutArray_188,
      S=>F_189, Cout=>CoutArray_189);
   forrow_11_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_175, Cin=>CoutArray_189,
      S=>F_190, Cout=>CoutArray_190);
   forrow_11_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_11_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_175, Cin=>
      CoutArray_190, S=>F_191, Cout=>CoutArray_191);
   forrow_12_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_177, Cin=>F_1024, S=>
      Product(12), Cout=>CoutArray_192);
   forrow_12_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_178, Cin=>CoutArray_192,
      S=>F_193, Cout=>CoutArray_193);
   forrow_12_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_179, Cin=>CoutArray_193,
      S=>F_194, Cout=>CoutArray_194);
   forrow_12_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_180, Cin=>CoutArray_194,
      S=>F_195, Cout=>CoutArray_195);
   forrow_12_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_181, Cin=>CoutArray_195,
      S=>F_196, Cout=>CoutArray_196);
   forrow_12_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_182, Cin=>CoutArray_196,
      S=>F_197, Cout=>CoutArray_197);
   forrow_12_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_183, Cin=>CoutArray_197,
      S=>F_198, Cout=>CoutArray_198);
   forrow_12_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_184, Cin=>CoutArray_198,
      S=>F_199, Cout=>CoutArray_199);
   forrow_12_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_185, Cin=>CoutArray_199,
      S=>F_200, Cout=>CoutArray_200);
   forrow_12_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_186, Cin=>CoutArray_200,
      S=>F_201, Cout=>CoutArray_201);
   forrow_12_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_187, Cin=>CoutArray_201,
      S=>F_202, Cout=>CoutArray_202);
   forrow_12_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_188, Cin=>CoutArray_202,
      S=>F_203, Cout=>CoutArray_203);
   forrow_12_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_189, Cin=>CoutArray_203,
      S=>F_204, Cout=>CoutArray_204);
   forrow_12_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_190, Cin=>CoutArray_204,
      S=>F_205, Cout=>CoutArray_205);
   forrow_12_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_191, Cin=>CoutArray_205,
      S=>F_206, Cout=>CoutArray_206);
   forrow_12_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_12_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_191, Cin=>
      CoutArray_206, S=>F_207, Cout=>CoutArray_207);
   forrow_13_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_193, Cin=>F_1024, S=>
      Product(13), Cout=>CoutArray_208);
   forrow_13_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_194, Cin=>CoutArray_208,
      S=>F_209, Cout=>CoutArray_209);
   forrow_13_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_195, Cin=>CoutArray_209,
      S=>F_210, Cout=>CoutArray_210);
   forrow_13_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_196, Cin=>CoutArray_210,
      S=>F_211, Cout=>CoutArray_211);
   forrow_13_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_197, Cin=>CoutArray_211,
      S=>F_212, Cout=>CoutArray_212);
   forrow_13_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_198, Cin=>CoutArray_212,
      S=>F_213, Cout=>CoutArray_213);
   forrow_13_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_199, Cin=>CoutArray_213,
      S=>F_214, Cout=>CoutArray_214);
   forrow_13_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_200, Cin=>CoutArray_214,
      S=>F_215, Cout=>CoutArray_215);
   forrow_13_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_201, Cin=>CoutArray_215,
      S=>F_216, Cout=>CoutArray_216);
   forrow_13_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_202, Cin=>CoutArray_216,
      S=>F_217, Cout=>CoutArray_217);
   forrow_13_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_203, Cin=>CoutArray_217,
      S=>F_218, Cout=>CoutArray_218);
   forrow_13_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_204, Cin=>CoutArray_218,
      S=>F_219, Cout=>CoutArray_219);
   forrow_13_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_205, Cin=>CoutArray_219,
      S=>F_220, Cout=>CoutArray_220);
   forrow_13_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_206, Cin=>CoutArray_220,
      S=>F_221, Cout=>CoutArray_221);
   forrow_13_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_207, Cin=>CoutArray_221,
      S=>F_222, Cout=>CoutArray_222);
   forrow_13_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_13_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_207, Cin=>
      CoutArray_222, S=>F_223, Cout=>CoutArray_223);
   forrow_14_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_209, Cin=>F_1024, S=>
      Product(14), Cout=>CoutArray_224);
   forrow_14_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_210, Cin=>CoutArray_224,
      S=>F_225, Cout=>CoutArray_225);
   forrow_14_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_211, Cin=>CoutArray_225,
      S=>F_226, Cout=>CoutArray_226);
   forrow_14_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_212, Cin=>CoutArray_226,
      S=>F_227, Cout=>CoutArray_227);
   forrow_14_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_213, Cin=>CoutArray_227,
      S=>F_228, Cout=>CoutArray_228);
   forrow_14_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_214, Cin=>CoutArray_228,
      S=>F_229, Cout=>CoutArray_229);
   forrow_14_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_215, Cin=>CoutArray_229,
      S=>F_230, Cout=>CoutArray_230);
   forrow_14_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_216, Cin=>CoutArray_230,
      S=>F_231, Cout=>CoutArray_231);
   forrow_14_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_217, Cin=>CoutArray_231,
      S=>F_232, Cout=>CoutArray_232);
   forrow_14_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_218, Cin=>CoutArray_232,
      S=>F_233, Cout=>CoutArray_233);
   forrow_14_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_219, Cin=>CoutArray_233,
      S=>F_234, Cout=>CoutArray_234);
   forrow_14_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_220, Cin=>CoutArray_234,
      S=>F_235, Cout=>CoutArray_235);
   forrow_14_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_221, Cin=>CoutArray_235,
      S=>F_236, Cout=>CoutArray_236);
   forrow_14_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_222, Cin=>CoutArray_236,
      S=>F_237, Cout=>CoutArray_237);
   forrow_14_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_223, Cin=>CoutArray_237,
      S=>F_238, Cout=>CoutArray_238);
   forrow_14_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_14_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_223, Cin=>
      CoutArray_238, S=>F_239, Cout=>CoutArray_239);
   forrow_15_ifn0_forcol_0_GEN0_ANDADD0_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_0_GEN0_ANDADD0_F, B=>F_225, Cin=>F_1024, S=>
      Product(15), Cout=>CoutArray_240);
   forrow_15_ifn0_forcol_1_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_1_GENX_ANDADDX_F, B=>F_226, Cin=>CoutArray_240,
      S=>Product(16), Cout=>CoutArray_241);
   forrow_15_ifn0_forcol_2_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_2_GENX_ANDADDX_F, B=>F_227, Cin=>CoutArray_241,
      S=>Product(17), Cout=>CoutArray_242);
   forrow_15_ifn0_forcol_3_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_3_GENX_ANDADDX_F, B=>F_228, Cin=>CoutArray_242,
      S=>Product(18), Cout=>CoutArray_243);
   forrow_15_ifn0_forcol_4_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_4_GENX_ANDADDX_F, B=>F_229, Cin=>CoutArray_243,
      S=>Product(19), Cout=>CoutArray_244);
   forrow_15_ifn0_forcol_5_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_5_GENX_ANDADDX_F, B=>F_230, Cin=>CoutArray_244,
      S=>Product(20), Cout=>CoutArray_245);
   forrow_15_ifn0_forcol_6_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_6_GENX_ANDADDX_F, B=>F_231, Cin=>CoutArray_245,
      S=>Product(21), Cout=>CoutArray_246);
   forrow_15_ifn0_forcol_7_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_7_GENX_ANDADDX_F, B=>F_232, Cin=>CoutArray_246,
      S=>Product(22), Cout=>CoutArray_247);
   forrow_15_ifn0_forcol_8_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_8_GENX_ANDADDX_F, B=>F_233, Cin=>CoutArray_247,
      S=>Product(23), Cout=>CoutArray_248);
   forrow_15_ifn0_forcol_9_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_9_GENX_ANDADDX_F, B=>F_234, Cin=>CoutArray_248,
      S=>Product(24), Cout=>CoutArray_249);
   forrow_15_ifn0_forcol_10_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_10_GENX_ANDADDX_F, B=>F_235, Cin=>CoutArray_249,
      S=>Product(25), Cout=>CoutArray_250);
   forrow_15_ifn0_forcol_11_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_11_GENX_ANDADDX_F, B=>F_236, Cin=>CoutArray_250,
      S=>Product(26), Cout=>CoutArray_251);
   forrow_15_ifn0_forcol_12_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_12_GENX_ANDADDX_F, B=>F_237, Cin=>CoutArray_251,
      S=>Product(27), Cout=>CoutArray_252);
   forrow_15_ifn0_forcol_13_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_13_GENX_ANDADDX_F, B=>F_238, Cin=>CoutArray_252,
      S=>Product(28), Cout=>CoutArray_253);
   forrow_15_ifn0_forcol_14_GENX_ANDADDX_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_14_GENX_ANDADDX_F, B=>F_239, Cin=>CoutArray_253,
      S=>Product(29), Cout=>CoutArray_254);
   forrow_15_ifn0_forcol_15_GENN_ANDADDN_FA : FA_1bit port map ( A=>
      forrow_15_ifn0_forcol_15_GENN_ANDADDN_F, B=>CoutArray_239, Cin=>
      CoutArray_254, S=>Product(30), Cout=>Product(31));
   ix1511 : fake_gnd port map ( Y=>F_1024);
   ix1 : and02 port map ( Y=>forrow_15_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(15), A1=>B(15));
   ix3 : and02 port map ( Y=>forrow_15_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(14));
   ix5 : and02 port map ( Y=>forrow_15_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(13));
   ix7 : and02 port map ( Y=>forrow_15_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(12));
   ix9 : and02 port map ( Y=>forrow_15_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(11));
   ix11 : and02 port map ( Y=>forrow_15_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(10));
   ix13 : and02 port map ( Y=>forrow_15_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(9));
   ix15 : and02 port map ( Y=>forrow_15_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(8));
   ix17 : and02 port map ( Y=>forrow_15_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(7));
   ix19 : and02 port map ( Y=>forrow_15_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(6));
   ix21 : and02 port map ( Y=>forrow_15_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(5));
   ix23 : and02 port map ( Y=>forrow_15_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(4));
   ix25 : and02 port map ( Y=>forrow_15_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(3));
   ix27 : and02 port map ( Y=>forrow_15_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(2));
   ix29 : and02 port map ( Y=>forrow_15_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(15), A1=>B(1));
   ix31 : and02 port map ( Y=>forrow_15_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(15), A1=>B(0));
   ix33 : and02 port map ( Y=>forrow_14_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(14), A1=>B(15));
   ix35 : and02 port map ( Y=>forrow_14_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(14));
   ix37 : and02 port map ( Y=>forrow_14_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(13));
   ix39 : and02 port map ( Y=>forrow_14_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(12));
   ix41 : and02 port map ( Y=>forrow_14_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(11));
   ix43 : and02 port map ( Y=>forrow_14_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(10));
   ix45 : and02 port map ( Y=>forrow_14_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(9));
   ix47 : and02 port map ( Y=>forrow_14_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(8));
   ix49 : and02 port map ( Y=>forrow_14_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(7));
   ix51 : and02 port map ( Y=>forrow_14_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(6));
   ix53 : and02 port map ( Y=>forrow_14_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(5));
   ix55 : and02 port map ( Y=>forrow_14_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(4));
   ix57 : and02 port map ( Y=>forrow_14_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(3));
   ix59 : and02 port map ( Y=>forrow_14_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(2));
   ix61 : and02 port map ( Y=>forrow_14_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(14), A1=>B(1));
   ix63 : and02 port map ( Y=>forrow_14_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(14), A1=>B(0));
   ix65 : and02 port map ( Y=>forrow_13_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(13), A1=>B(15));
   ix67 : and02 port map ( Y=>forrow_13_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(14));
   ix69 : and02 port map ( Y=>forrow_13_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(13));
   ix71 : and02 port map ( Y=>forrow_13_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(12));
   ix73 : and02 port map ( Y=>forrow_13_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(11));
   ix75 : and02 port map ( Y=>forrow_13_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(10));
   ix77 : and02 port map ( Y=>forrow_13_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(9));
   ix79 : and02 port map ( Y=>forrow_13_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(8));
   ix81 : and02 port map ( Y=>forrow_13_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(7));
   ix83 : and02 port map ( Y=>forrow_13_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(6));
   ix85 : and02 port map ( Y=>forrow_13_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(5));
   ix87 : and02 port map ( Y=>forrow_13_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(4));
   ix89 : and02 port map ( Y=>forrow_13_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(3));
   ix91 : and02 port map ( Y=>forrow_13_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(2));
   ix93 : and02 port map ( Y=>forrow_13_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(13), A1=>B(1));
   ix95 : and02 port map ( Y=>forrow_13_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(13), A1=>B(0));
   ix97 : and02 port map ( Y=>forrow_12_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(12), A1=>B(15));
   ix99 : and02 port map ( Y=>forrow_12_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(14));
   ix101 : and02 port map ( Y=>forrow_12_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(13));
   ix103 : and02 port map ( Y=>forrow_12_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(12));
   ix105 : and02 port map ( Y=>forrow_12_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(11));
   ix107 : and02 port map ( Y=>forrow_12_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(10));
   ix109 : and02 port map ( Y=>forrow_12_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(9));
   ix111 : and02 port map ( Y=>forrow_12_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(8));
   ix113 : and02 port map ( Y=>forrow_12_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(7));
   ix115 : and02 port map ( Y=>forrow_12_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(6));
   ix117 : and02 port map ( Y=>forrow_12_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(5));
   ix119 : and02 port map ( Y=>forrow_12_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(4));
   ix121 : and02 port map ( Y=>forrow_12_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(3));
   ix123 : and02 port map ( Y=>forrow_12_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(2));
   ix125 : and02 port map ( Y=>forrow_12_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(12), A1=>B(1));
   ix127 : and02 port map ( Y=>forrow_12_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(12), A1=>B(0));
   ix129 : and02 port map ( Y=>forrow_11_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(11), A1=>B(15));
   ix131 : and02 port map ( Y=>forrow_11_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(14));
   ix133 : and02 port map ( Y=>forrow_11_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(13));
   ix135 : and02 port map ( Y=>forrow_11_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(12));
   ix137 : and02 port map ( Y=>forrow_11_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(11));
   ix139 : and02 port map ( Y=>forrow_11_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(10));
   ix141 : and02 port map ( Y=>forrow_11_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(9));
   ix143 : and02 port map ( Y=>forrow_11_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(8));
   ix145 : and02 port map ( Y=>forrow_11_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(7));
   ix147 : and02 port map ( Y=>forrow_11_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(6));
   ix149 : and02 port map ( Y=>forrow_11_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(5));
   ix151 : and02 port map ( Y=>forrow_11_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(4));
   ix153 : and02 port map ( Y=>forrow_11_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(3));
   ix155 : and02 port map ( Y=>forrow_11_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(2));
   ix157 : and02 port map ( Y=>forrow_11_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(11), A1=>B(1));
   ix159 : and02 port map ( Y=>forrow_11_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(11), A1=>B(0));
   ix161 : and02 port map ( Y=>forrow_10_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(10), A1=>B(15));
   ix163 : and02 port map ( Y=>forrow_10_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(14));
   ix165 : and02 port map ( Y=>forrow_10_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(13));
   ix167 : and02 port map ( Y=>forrow_10_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(12));
   ix169 : and02 port map ( Y=>forrow_10_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(11));
   ix171 : and02 port map ( Y=>forrow_10_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(10));
   ix173 : and02 port map ( Y=>forrow_10_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(9));
   ix175 : and02 port map ( Y=>forrow_10_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(8));
   ix177 : and02 port map ( Y=>forrow_10_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(7));
   ix179 : and02 port map ( Y=>forrow_10_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(6));
   ix181 : and02 port map ( Y=>forrow_10_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(5));
   ix183 : and02 port map ( Y=>forrow_10_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(4));
   ix185 : and02 port map ( Y=>forrow_10_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(3));
   ix187 : and02 port map ( Y=>forrow_10_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(2));
   ix189 : and02 port map ( Y=>forrow_10_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(10), A1=>B(1));
   ix191 : and02 port map ( Y=>forrow_10_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(10), A1=>B(0));
   ix193 : and02 port map ( Y=>forrow_9_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(9), A1=>B(15));
   ix195 : and02 port map ( Y=>forrow_9_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(14));
   ix197 : and02 port map ( Y=>forrow_9_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(13));
   ix199 : and02 port map ( Y=>forrow_9_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(12));
   ix201 : and02 port map ( Y=>forrow_9_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(11));
   ix203 : and02 port map ( Y=>forrow_9_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(10));
   ix205 : and02 port map ( Y=>forrow_9_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(9));
   ix207 : and02 port map ( Y=>forrow_9_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(8));
   ix209 : and02 port map ( Y=>forrow_9_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(7));
   ix211 : and02 port map ( Y=>forrow_9_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(6));
   ix213 : and02 port map ( Y=>forrow_9_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(5));
   ix215 : and02 port map ( Y=>forrow_9_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(4));
   ix217 : and02 port map ( Y=>forrow_9_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(3));
   ix219 : and02 port map ( Y=>forrow_9_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(2));
   ix221 : and02 port map ( Y=>forrow_9_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(9), A1=>B(1));
   ix223 : and02 port map ( Y=>forrow_9_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(9), A1=>B(0));
   ix225 : and02 port map ( Y=>forrow_8_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(8), A1=>B(15));
   ix227 : and02 port map ( Y=>forrow_8_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(14));
   ix229 : and02 port map ( Y=>forrow_8_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(13));
   ix231 : and02 port map ( Y=>forrow_8_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(12));
   ix233 : and02 port map ( Y=>forrow_8_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(11));
   ix235 : and02 port map ( Y=>forrow_8_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(10));
   ix237 : and02 port map ( Y=>forrow_8_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(9));
   ix239 : and02 port map ( Y=>forrow_8_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(8));
   ix241 : and02 port map ( Y=>forrow_8_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(7));
   ix243 : and02 port map ( Y=>forrow_8_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(6));
   ix245 : and02 port map ( Y=>forrow_8_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(5));
   ix247 : and02 port map ( Y=>forrow_8_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(4));
   ix249 : and02 port map ( Y=>forrow_8_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(3));
   ix251 : and02 port map ( Y=>forrow_8_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(2));
   ix253 : and02 port map ( Y=>forrow_8_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(8), A1=>B(1));
   ix255 : and02 port map ( Y=>forrow_8_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(8), A1=>B(0));
   ix257 : and02 port map ( Y=>forrow_7_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(7), A1=>B(15));
   ix259 : and02 port map ( Y=>forrow_7_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(14));
   ix261 : and02 port map ( Y=>forrow_7_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(13));
   ix263 : and02 port map ( Y=>forrow_7_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(12));
   ix265 : and02 port map ( Y=>forrow_7_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(11));
   ix267 : and02 port map ( Y=>forrow_7_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(10));
   ix269 : and02 port map ( Y=>forrow_7_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(9));
   ix271 : and02 port map ( Y=>forrow_7_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(8));
   ix273 : and02 port map ( Y=>forrow_7_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(7));
   ix275 : and02 port map ( Y=>forrow_7_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(6));
   ix277 : and02 port map ( Y=>forrow_7_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(5));
   ix279 : and02 port map ( Y=>forrow_7_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(4));
   ix281 : and02 port map ( Y=>forrow_7_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(3));
   ix283 : and02 port map ( Y=>forrow_7_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(2));
   ix285 : and02 port map ( Y=>forrow_7_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(7), A1=>B(1));
   ix287 : and02 port map ( Y=>forrow_7_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(7), A1=>B(0));
   ix289 : and02 port map ( Y=>forrow_6_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(6), A1=>B(15));
   ix291 : and02 port map ( Y=>forrow_6_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(14));
   ix293 : and02 port map ( Y=>forrow_6_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(13));
   ix295 : and02 port map ( Y=>forrow_6_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(12));
   ix297 : and02 port map ( Y=>forrow_6_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(11));
   ix299 : and02 port map ( Y=>forrow_6_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(10));
   ix301 : and02 port map ( Y=>forrow_6_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(9));
   ix303 : and02 port map ( Y=>forrow_6_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(8));
   ix305 : and02 port map ( Y=>forrow_6_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(7));
   ix307 : and02 port map ( Y=>forrow_6_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(6));
   ix309 : and02 port map ( Y=>forrow_6_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(5));
   ix311 : and02 port map ( Y=>forrow_6_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(4));
   ix313 : and02 port map ( Y=>forrow_6_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(3));
   ix315 : and02 port map ( Y=>forrow_6_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(2));
   ix317 : and02 port map ( Y=>forrow_6_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(6), A1=>B(1));
   ix319 : and02 port map ( Y=>forrow_6_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(6), A1=>B(0));
   ix321 : and02 port map ( Y=>forrow_5_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(5), A1=>B(15));
   ix323 : and02 port map ( Y=>forrow_5_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(14));
   ix325 : and02 port map ( Y=>forrow_5_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(13));
   ix327 : and02 port map ( Y=>forrow_5_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(12));
   ix329 : and02 port map ( Y=>forrow_5_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(11));
   ix331 : and02 port map ( Y=>forrow_5_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(10));
   ix333 : and02 port map ( Y=>forrow_5_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(9));
   ix335 : and02 port map ( Y=>forrow_5_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(8));
   ix337 : and02 port map ( Y=>forrow_5_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(7));
   ix339 : and02 port map ( Y=>forrow_5_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(6));
   ix341 : and02 port map ( Y=>forrow_5_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(5));
   ix343 : and02 port map ( Y=>forrow_5_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(4));
   ix345 : and02 port map ( Y=>forrow_5_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(3));
   ix347 : and02 port map ( Y=>forrow_5_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(2));
   ix349 : and02 port map ( Y=>forrow_5_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(5), A1=>B(1));
   ix351 : and02 port map ( Y=>forrow_5_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(5), A1=>B(0));
   ix353 : and02 port map ( Y=>forrow_4_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(4), A1=>B(15));
   ix355 : and02 port map ( Y=>forrow_4_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(14));
   ix357 : and02 port map ( Y=>forrow_4_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(13));
   ix359 : and02 port map ( Y=>forrow_4_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(12));
   ix361 : and02 port map ( Y=>forrow_4_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(11));
   ix363 : and02 port map ( Y=>forrow_4_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(10));
   ix365 : and02 port map ( Y=>forrow_4_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(9));
   ix367 : and02 port map ( Y=>forrow_4_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(8));
   ix369 : and02 port map ( Y=>forrow_4_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(7));
   ix371 : and02 port map ( Y=>forrow_4_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(6));
   ix373 : and02 port map ( Y=>forrow_4_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(5));
   ix375 : and02 port map ( Y=>forrow_4_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(4));
   ix377 : and02 port map ( Y=>forrow_4_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(3));
   ix379 : and02 port map ( Y=>forrow_4_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(2));
   ix381 : and02 port map ( Y=>forrow_4_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(4), A1=>B(1));
   ix383 : and02 port map ( Y=>forrow_4_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(4), A1=>B(0));
   ix385 : and02 port map ( Y=>forrow_3_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(3), A1=>B(15));
   ix387 : and02 port map ( Y=>forrow_3_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(14));
   ix389 : and02 port map ( Y=>forrow_3_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(13));
   ix391 : and02 port map ( Y=>forrow_3_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(12));
   ix393 : and02 port map ( Y=>forrow_3_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(11));
   ix395 : and02 port map ( Y=>forrow_3_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(10));
   ix397 : and02 port map ( Y=>forrow_3_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(9));
   ix399 : and02 port map ( Y=>forrow_3_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(8));
   ix401 : and02 port map ( Y=>forrow_3_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(7));
   ix403 : and02 port map ( Y=>forrow_3_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(6));
   ix405 : and02 port map ( Y=>forrow_3_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(5));
   ix407 : and02 port map ( Y=>forrow_3_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(4));
   ix409 : and02 port map ( Y=>forrow_3_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(3));
   ix411 : and02 port map ( Y=>forrow_3_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(2));
   ix413 : and02 port map ( Y=>forrow_3_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(3), A1=>B(1));
   ix415 : and02 port map ( Y=>forrow_3_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(3), A1=>B(0));
   ix417 : and02 port map ( Y=>forrow_2_ifn0_forcol_15_GENN_ANDADDN_F, A0=>
      A(2), A1=>B(15));
   ix419 : and02 port map ( Y=>forrow_2_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(14));
   ix421 : and02 port map ( Y=>forrow_2_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(13));
   ix423 : and02 port map ( Y=>forrow_2_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(12));
   ix425 : and02 port map ( Y=>forrow_2_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(11));
   ix427 : and02 port map ( Y=>forrow_2_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(10));
   ix429 : and02 port map ( Y=>forrow_2_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(9));
   ix431 : and02 port map ( Y=>forrow_2_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(8));
   ix433 : and02 port map ( Y=>forrow_2_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(7));
   ix435 : and02 port map ( Y=>forrow_2_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(6));
   ix437 : and02 port map ( Y=>forrow_2_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(5));
   ix439 : and02 port map ( Y=>forrow_2_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(4));
   ix441 : and02 port map ( Y=>forrow_2_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(3));
   ix443 : and02 port map ( Y=>forrow_2_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(2));
   ix445 : and02 port map ( Y=>forrow_2_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(2), A1=>B(1));
   ix447 : and02 port map ( Y=>forrow_2_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(2), A1=>B(0));
   ix449 : and02 port map ( Y=>forrow_1_ifn0_forcol_15_GEN1N_ANDADD1N_F, A0
      =>A(1), A1=>B(15));
   ix451 : and02 port map ( Y=>forrow_1_ifn0_forcol_14_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(14));
   ix453 : and02 port map ( Y=>forrow_1_ifn0_forcol_13_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(13));
   ix455 : and02 port map ( Y=>forrow_1_ifn0_forcol_12_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(12));
   ix457 : and02 port map ( Y=>forrow_1_ifn0_forcol_11_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(11));
   ix459 : and02 port map ( Y=>forrow_1_ifn0_forcol_10_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(10));
   ix461 : and02 port map ( Y=>forrow_1_ifn0_forcol_9_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(9));
   ix463 : and02 port map ( Y=>forrow_1_ifn0_forcol_8_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(8));
   ix465 : and02 port map ( Y=>forrow_1_ifn0_forcol_7_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(7));
   ix467 : and02 port map ( Y=>forrow_1_ifn0_forcol_6_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(6));
   ix469 : and02 port map ( Y=>forrow_1_ifn0_forcol_5_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(5));
   ix471 : and02 port map ( Y=>forrow_1_ifn0_forcol_4_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(4));
   ix473 : and02 port map ( Y=>forrow_1_ifn0_forcol_3_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(3));
   ix475 : and02 port map ( Y=>forrow_1_ifn0_forcol_2_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(2));
   ix477 : and02 port map ( Y=>forrow_1_ifn0_forcol_1_GENX_ANDADDX_F, A0=>
      A(1), A1=>B(1));
   ix479 : and02 port map ( Y=>forrow_1_ifn0_forcol_0_GEN0_ANDADD0_F, A0=>
      A(1), A1=>B(0));
   ix509 : and02 port map ( Y=>F_1, A0=>B(1), A1=>A(0));
   ix507 : and02 port map ( Y=>F_2, A0=>B(2), A1=>A(0));
   ix505 : and02 port map ( Y=>F_3, A0=>B(3), A1=>A(0));
   ix503 : and02 port map ( Y=>F_4, A0=>B(4), A1=>A(0));
   ix501 : and02 port map ( Y=>F_5, A0=>B(5), A1=>A(0));
   ix499 : and02 port map ( Y=>F_6, A0=>B(6), A1=>A(0));
   ix497 : and02 port map ( Y=>F_7, A0=>B(7), A1=>A(0));
   ix495 : and02 port map ( Y=>F_8, A0=>B(8), A1=>A(0));
   ix493 : and02 port map ( Y=>F_9, A0=>B(9), A1=>A(0));
   ix491 : and02 port map ( Y=>F_10, A0=>B(10), A1=>A(0));
   ix489 : and02 port map ( Y=>F_11, A0=>B(11), A1=>A(0));
   ix487 : and02 port map ( Y=>F_12, A0=>B(12), A1=>A(0));
   ix485 : and02 port map ( Y=>F_13, A0=>B(13), A1=>A(0));
   ix483 : and02 port map ( Y=>F_14, A0=>B(14), A1=>A(0));
   ix481 : and02 port map ( Y=>F_15, A0=>B(15), A1=>A(0));
   ix511 : and02 port map ( Y=>Product(0), A0=>B(0), A1=>A(0));
end Behavioral ;

