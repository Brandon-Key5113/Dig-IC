* Example circuit file for simulating PEX

.OPTION DOTNODE
.HIER /

.INCLUDE "/home/bxk5113/Pyxis_SPT_HEP/ic_projects/Pyxis_SPT/digicdesign/ProjectWrapper/ProjectWrapper.cal/ProjectWrapper.pex.netlist"

.LIB /home/bxk5113/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT

* - Instantiate your parasitic netlist and add the load capacitor
** FORMAT :
* XLAYOUT [all inputs as listed by the ".subckt" line in the included netlist, in the order that they appear there] [name of the subcircuit as listed in the included netlist]
XLAYOUT COMPLETE PASS REGOUT[31] REGOUT[30] REGOUT[29] REGOUT[28] REGOUT[27] REGOUT[26] REGOUT[25] REGOUT[24] REGOUT[23] REGOUT[22] REGOUT[21] REGOUT[20] REGOUT[19] REGOUT[18] REGOUT[17] REGOUT[16] REGOUT[15] REGOUT[14] REGOUT[13] REGOUT[12] REGOUT[11] REGOUT[10] REGOUT[9] REGOUT[8] REGOUT[7] REGOUT[6] REGOUT[5] REGOUT[4] REGOUT[3] REGOUT[2] REGOUT[1] REGOUT[0] A[15] A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CLK RESET STARTTEST WE ProjectWrapper

* Output Capactitance
C_REGOUT[31] REGOUT[31] 0 120f
C_REGOUT[30] REGOUT[30] 0 120f
C_REGOUT[29] REGOUT[29] 0 120f
C_REGOUT[28] REGOUT[28] 0 120f
C_REGOUT[27] REGOUT[27] 0 120f
C_REGOUT[26] REGOUT[26] 0 120f
C_REGOUT[25] REGOUT[25] 0 120f
C_REGOUT[24] REGOUT[24] 0 120f
C_REGOUT[23] REGOUT[23] 0 120f
C_REGOUT[22] REGOUT[22] 0 120f
C_REGOUT[21] REGOUT[21] 0 120f
C_REGOUT[20] REGOUT[20] 0 120f
C_REGOUT[19] REGOUT[19] 0 120f
C_REGOUT[18] REGOUT[18] 0 120f
C_REGOUT[17] REGOUT[17] 0 120f
C_REGOUT[16] REGOUT[16] 0 120f
C_REGOUT[15] REGOUT[15] 0 120f
C_REGOUT[14] REGOUT[14] 0 120f
C_REGOUT[13] REGOUT[13] 0 120f
C_REGOUT[12] REGOUT[12] 0 120f
C_REGOUT[11] REGOUT[11] 0 120f
C_REGOUT[10] REGOUT[10] 0 120f
C_REGOUT[9] REGOUT[9] 0 120f
C_REGOUT[8] REGOUT[8] 0 120f
C_REGOUT[7] REGOUT[7] 0 120f
C_REGOUT[6] REGOUT[6] 0 120f
C_REGOUT[5] REGOUT[5] 0 120f
C_REGOUT[4] REGOUT[4] 0 120f
C_REGOUT[3] REGOUT[3] 0 120f
C_REGOUT[2] REGOUT[2] 0 120f
C_REGOUT[1] REGOUT[1] 0 120f
C_REGOUT[0] REGOUT[0] 0 120f


* - Analysis Setup - DC sweep
* FORMAT : .DC [name] [low] [high] [step]
*.DC VFORCE__A 0 1.2 0.01

* - Analysis Setup - Trans
* FORMAT : .TRAN [start time] [end time] [time step]
.TRAN 0 2000n 0.05n

* --- Forces
* FORMAT -- PULSE : [name] [port] [reference (0 means ground)] PULSE [low] [high] [delay] [fall time] [rise time] [pulse width] [period]
*
* FORMAT -- DC    : [name] [port] [reference (0 means ground)] DC [voltage]
*

VFORCE__VDD VDD 0 DC 1.08
VFORCE__VSS VSS 0 DC 0

VFORCE__CLK CLK 0 PULSE (0 1.08 25n 0.1n 0.1n 25n 50n)

VFORCE__RESET RESET 0 pwl (120n 1.08 120.1n 0 )
VFORCE__WE WE 0 DC 1.08

.SIGBUS A[15:0] VHI=1.08 VLO=0 TRISE=0.1n TFALL=0.1n TDELAY=210n THOLD=200n BASE=HEXA PATTERN 0002 0003 P
.SIGBUS B[15:0] VHI=1.08 VLO=0 TRISE=0.1n TFALL=0.1n TDELAY=210n THOLD=200n BASE=HEXA PATTERN 0003 0004 P


* --- Waveform Outputs
.PLOT TRAN V(COMPLETE)
.PLOT TRAN V(PASS)
.PLOT TRAN V(REGOUT[31])
.PLOT TRAN V(REGOUT[30])
.PLOT TRAN V(REGOUT[29])
.PLOT TRAN V(REGOUT[28])
.PLOT TRAN V(REGOUT[27])
.PLOT TRAN V(REGOUT[26])
.PLOT TRAN V(REGOUT[25])
.PLOT TRAN V(REGOUT[24])
.PLOT TRAN V(REGOUT[23])
.PLOT TRAN V(REGOUT[22])
.PLOT TRAN V(REGOUT[21])
.PLOT TRAN V(REGOUT[20])
.PLOT TRAN V(REGOUT[19])
.PLOT TRAN V(REGOUT[18])
.PLOT TRAN V(REGOUT[17])
.PLOT TRAN V(REGOUT[16])
.PLOT TRAN V(REGOUT[15])
.PLOT TRAN V(REGOUT[14])
.PLOT TRAN V(REGOUT[13])
.PLOT TRAN V(REGOUT[12])
.PLOT TRAN V(REGOUT[11])
.PLOT TRAN V(REGOUT[10])
.PLOT TRAN V(REGOUT[9])
.PLOT TRAN V(REGOUT[8])
.PLOT TRAN V(REGOUT[7])
.PLOT TRAN V(REGOUT[6])
.PLOT TRAN V(REGOUT[5])
.PLOT TRAN V(REGOUT[4])
.PLOT TRAN V(REGOUT[3])
.PLOT TRAN V(REGOUT[2])
.PLOT TRAN V(REGOUT[1])
.PLOT TRAN V(REGOUT[0])
.PLOT TRAN V(A[15])
.PLOT TRAN V(A[14])
.PLOT TRAN V(A[13])
.PLOT TRAN V(A[12])
.PLOT TRAN V(A[11])
.PLOT TRAN V(A[10])
.PLOT TRAN V(A[9])
.PLOT TRAN V(A[8])
.PLOT TRAN V(A[7])
.PLOT TRAN V(A[6])
.PLOT TRAN V(A[5])
.PLOT TRAN V(A[4])
.PLOT TRAN V(A[3])
.PLOT TRAN V(A[2])
.PLOT TRAN V(A[1])
.PLOT TRAN V(A[0])
.PLOT TRAN V(B[15])
.PLOT TRAN V(B[14])
.PLOT TRAN V(B[13])
.PLOT TRAN V(B[12])
.PLOT TRAN V(B[11])
.PLOT TRAN V(B[10])
.PLOT TRAN V(B[9])
.PLOT TRAN V(B[8])
.PLOT TRAN V(B[7])
.PLOT TRAN V(B[6])
.PLOT TRAN V(B[5])
.PLOT TRAN V(B[4])
.PLOT TRAN V(B[3])
.PLOT TRAN V(B[2])
.PLOT TRAN V(B[1])
.PLOT TRAN V(B[0])
.PLOT TRAN V(CLK)
.PLOT TRAN V(RESET)
.PLOT TRAN V(STARTTEST)
.PLOT TRAN V(WE)


* --- Params
.TEMP 125

* --- Power Measurement
.measure tran static_pwr AVG power from=90ns to=160ns
.measure tran inst_pwr MAX power from=90ns to=160ns

