* Component: $PYXIS_SPT/digicdesign/mirroradder Viewpoint: default

.INCLUDE "$PYXIS_SPT/digicdesign/mirroradder/default/netlist.spi"
.INCLUDE "$GENERIC13/models/include_all"
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - DCOP
.OPTION PROBEOP2
.OP

* - Analysis Setup - Trans
.TRAN 0 160n 0n

* --- Forces
VFORCE__A A GROUND PULSE (0 1.08 20n .1n .1n 20n 40n)
VFORCE__B B GROUND PULSE (0 1.08 40n .1n .1n 40n 80n)
VFORCE__Cin CIN GROUND PULSE (0 1.08 80n .1n .1n 80n 160n)
VFORCE__Vdd VDD GROUND DC 1.08

* --- Global Outputs
.PROBE V SG

* --- Params
.TEMP 125.0

* --- Libsetup
.LIB KEY=MOS "$GENERIC13/models/lib.eldo" TT
.LIB KEY=MOS_33 "$GENERIC13/models/lib.eldo" TT_33
.LIB KEY=MOS_lvt "$GENERIC13/models/lib.eldo" TT_lvt
.LIB KEY=MOS_hvt "$GENERIC13/models/lib.eldo" TT_hvt
.LIB KEY=BIP "$GENERIC13/models/lib.eldo" TT_BIP
.LIB KEY=BIP_NPN "$GENERIC13/models/lib.eldo" TT_BIP_NPN
.LIB KEY=RES "$GENERIC13/models/lib.eldo" TT_RES
