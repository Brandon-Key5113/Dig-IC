
-- 
-- Definition of  nBitAND_4Bit
-- 
--      Sun Nov  3 13:53:06 2019
--      
--      LeonardoSpectrum Level 3, 2008b.3
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity nBitAND_4Bit is
   port (
      A : IN std_logic_vector (15 DOWNTO 0) ;
      B : IN std_logic_vector (15 DOWNTO 0) ;
      Y : OUT std_logic_vector (15 DOWNTO 0)) ;
end nBitAND_4Bit ;

architecture Dataflow of nBitAND_4Bit is
begin
   ix1 : and02 port map ( Y=>Y(0), A0=>B(0), A1=>A(0));
   ix3 : and02 port map ( Y=>Y(1), A0=>B(1), A1=>A(1));
   ix5 : and02 port map ( Y=>Y(2), A0=>B(2), A1=>A(2));
   ix7 : and02 port map ( Y=>Y(3), A0=>B(3), A1=>A(3));
   ix9 : and02 port map ( Y=>Y(4), A0=>B(4), A1=>A(4));
   ix11 : and02 port map ( Y=>Y(5), A0=>B(5), A1=>A(5));
   ix13 : and02 port map ( Y=>Y(6), A0=>B(6), A1=>A(6));
   ix15 : and02 port map ( Y=>Y(7), A0=>B(7), A1=>A(7));
   ix17 : and02 port map ( Y=>Y(8), A0=>B(8), A1=>A(8));
   ix19 : and02 port map ( Y=>Y(9), A0=>B(9), A1=>A(9));
   ix21 : and02 port map ( Y=>Y(10), A0=>B(10), A1=>A(10));
   ix23 : and02 port map ( Y=>Y(11), A0=>B(11), A1=>A(11));
   ix25 : and02 port map ( Y=>Y(12), A0=>B(12), A1=>A(12));
   ix27 : and02 port map ( Y=>Y(13), A0=>B(13), A1=>A(13));
   ix29 : and02 port map ( Y=>Y(14), A0=>B(14), A1=>A(14));
   ix31 : and02 port map ( Y=>Y(15), A0=>B(15), A1=>A(15));
end Dataflow ;

