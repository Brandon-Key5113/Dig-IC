* SPICE NETLIST
***************************************

.SUBCKT mimcap_g13 plus minus
.ENDS
***************************************
.SUBCKT spiral_inductor_lvs pos neg
.ENDS
***************************************
.SUBCKT inv01 VSS VDD Y A
** N=4 EP=4 IP=0 FDC=2
M0 Y A VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=910 $Y=1820 $D=19
M1 Y A VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=910 $Y=5600 $D=25
.ENDS
***************************************
.SUBCKT or02 VSS VDD Y A1 A0
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=805 $Y=1330 $D=19
M1 VSS A0 6 VSS nmos L=1.4e-07 W=3.5e-07 $X=1365 $Y=1330 $D=19
M2 Y 6 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=1925 $Y=1330 $D=19
M3 7 A1 6 VDD pmos L=1.4e-07 W=1.19e-06 $X=910 $Y=5880 $D=25
M4 VDD A0 7 VDD pmos L=1.4e-07 W=1.19e-06 $X=1330 $Y=5880 $D=25
M5 Y 6 VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=1925 $Y=5880 $D=25
.ENDS
***************************************
.SUBCKT nand02 VSS Y VDD A1 A0
** N=6 EP=5 IP=0 FDC=4
M0 6 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=875 $Y=1190 $D=19
M1 Y A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=1295 $Y=1190 $D=19
M2 Y A1 VDD VDD pmos L=1.4e-07 W=1.05e-06 $X=875 $Y=6160 $D=25
M3 VDD A0 Y VDD pmos L=1.4e-07 W=1.05e-06 $X=1435 $Y=6160 $D=25
.ENDS
***************************************
.SUBCKT oai321 VDD Y VSS A0 A1 A2 B1 B0 C0
** N=14 EP=9 IP=0 FDC=12
M0 10 A0 Y VSS nmos L=1.4e-07 W=1.19e-06 $X=805 $Y=1295 $D=19
M1 Y A1 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=1365 $Y=1295 $D=19
M2 10 A2 Y VSS nmos L=1.4e-07 W=1.19e-06 $X=1925 $Y=1295 $D=19
M3 10 B1 11 VSS nmos L=1.4e-07 W=1.19e-06 $X=3045 $Y=1295 $D=19
M4 11 B0 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=3605 $Y=1295 $D=19
M5 VSS C0 11 VSS nmos L=1.4e-07 W=1.19e-06 $X=4165 $Y=1295 $D=19
M6 12 A0 VDD VDD pmos L=1.4e-07 W=3.15e-06 $X=1260 $Y=4060 $D=25
M7 13 A1 12 VDD pmos L=1.4e-07 W=3.15e-06 $X=1680 $Y=4060 $D=25
M8 Y A2 13 VDD pmos L=1.4e-07 W=3.15e-06 $X=2100 $Y=4060 $D=25
M9 14 B1 Y VDD pmos L=1.4e-07 W=2.24e-06 $X=2695 $Y=4970 $D=25
M10 VDD B0 14 VDD pmos L=1.4e-07 W=2.24e-06 $X=3115 $Y=4970 $D=25
M11 Y C0 VDD VDD pmos L=1.4e-07 W=1.26e-06 $X=3710 $Y=4970 $D=25
.ENDS
***************************************
.SUBCKT xor2 VSS VDD Y A1 A0
** N=10 EP=5 IP=0 FDC=12
M0 7 A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1330 $D=19
M1 VSS A1 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1225 $Y=1330 $D=19
M2 8 6 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=1785 $Y=1330 $D=19
M3 9 A1 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=2345 $Y=1330 $D=19
M4 8 A0 9 VSS nmos L=1.4e-07 W=7.7e-07 $X=2905 $Y=1330 $D=19
M5 Y 9 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=4025 $Y=1330 $D=19
M6 6 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=875 $Y=5880 $D=25
M7 VDD A1 6 VDD pmos L=1.4e-07 W=1.19e-06 $X=1435 $Y=5880 $D=25
M8 9 6 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1995 $Y=5880 $D=25
M9 10 A1 9 VDD pmos L=1.4e-07 W=2.24e-06 $X=2590 $Y=4830 $D=25
M10 VDD A0 10 VDD pmos L=1.4e-07 W=2.24e-06 $X=3010 $Y=4830 $D=25
M11 Y 9 VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=3605 $Y=4830 $D=25
.ENDS
***************************************
.SUBCKT nor03 Y VDD VSS A0 A1 A2
** N=8 EP=6 IP=0 FDC=6
M0 VSS A0 Y VSS nmos L=1.4e-07 W=4.2e-07 $X=875 $Y=1190 $D=19
M1 Y A1 VSS VSS nmos L=1.4e-07 W=4.2e-07 $X=1435 $Y=1190 $D=19
M2 VSS A2 Y VSS nmos L=1.4e-07 W=4.2e-07 $X=1995 $Y=1190 $D=19
M3 7 A0 VDD VDD pmos L=1.4e-07 W=1.68e-06 $X=875 $Y=5530 $D=25
M4 8 A1 7 VDD pmos L=1.4e-07 W=1.68e-06 $X=1295 $Y=5530 $D=25
M5 Y A2 8 VDD pmos L=1.4e-07 W=1.68e-06 $X=1715 $Y=5530 $D=25
.ENDS
***************************************
.SUBCKT aoi22 VSS VDD Y A1 A0 B0 B1
** N=10 EP=7 IP=0 FDC=8
M0 8 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=945 $Y=1190 $D=19
M1 Y A0 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=1365 $Y=1190 $D=19
M2 9 B0 Y VSS nmos L=1.4e-07 W=7.7e-07 $X=1925 $Y=1190 $D=19
M3 VSS B1 9 VSS nmos L=1.4e-07 W=7.7e-07 $X=2345 $Y=1190 $D=19
M4 VDD A1 10 VDD pmos L=1.4e-07 W=1.19e-06 $X=805 $Y=6020 $D=25
M5 10 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1365 $Y=6020 $D=25
M6 Y B0 10 VDD pmos L=1.4e-07 W=1.19e-06 $X=1925 $Y=6020 $D=25
M7 10 B1 Y VDD pmos L=1.4e-07 W=1.19e-06 $X=2485 $Y=6020 $D=25
.ENDS
***************************************
.SUBCKT nor02ii VSS VDD Y A1 A0
** N=7 EP=5 IP=0 FDC=6
M0 VSS A1 6 VSS nmos L=1.4e-07 W=3.5e-07 $X=805 $Y=1190 $D=19
M1 Y A0 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=1365 $Y=1190 $D=19
M2 VSS 6 Y VSS nmos L=1.4e-07 W=3.5e-07 $X=1925 $Y=1190 $D=19
M3 VDD A1 6 VDD pmos L=1.4e-07 W=7.7e-07 $X=805 $Y=6020 $D=25
M4 7 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1400 $Y=6020 $D=25
M5 Y 6 7 VDD pmos L=1.4e-07 W=1.19e-06 $X=1820 $Y=6020 $D=25
.ENDS
***************************************
.SUBCKT oai21 VSS Y VDD B0 A1 A0
** N=8 EP=6 IP=0 FDC=6
M0 7 B0 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1235 $D=19
M1 Y A1 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1365 $Y=1235 $D=19
M2 7 A0 Y VSS nmos L=1.4e-07 W=7.7e-07 $X=1925 $Y=1235 $D=19
M3 Y B0 VDD VDD pmos L=1.4e-07 W=1.05e-06 $X=910 $Y=5180 $D=25
M4 8 A1 Y VDD pmos L=1.4e-07 W=2.03e-06 $X=1505 $Y=5180 $D=25
M5 VDD A0 8 VDD pmos L=1.4e-07 W=2.03e-06 $X=1925 $Y=5180 $D=25
.ENDS
***************************************
.SUBCKT ao22 VSS VDD Y A1 B0 B1 A0
** N=11 EP=7 IP=0 FDC=10
M0 8 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=945 $Y=1190 $D=19
M1 9 A0 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=1365 $Y=1190 $D=19
M2 10 B0 9 VSS nmos L=1.4e-07 W=7.7e-07 $X=1925 $Y=1190 $D=19
M3 VSS B1 10 VSS nmos L=1.4e-07 W=7.7e-07 $X=2345 $Y=1190 $D=19
M4 Y 9 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=2940 $Y=1610 $D=19
M5 11 A1 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=805 $Y=6020 $D=25
M6 9 B0 11 VDD pmos L=1.4e-07 W=1.19e-06 $X=1365 $Y=6020 $D=25
M7 11 B1 9 VDD pmos L=1.4e-07 W=1.19e-06 $X=1925 $Y=6020 $D=25
M8 VDD A0 11 VDD pmos L=1.4e-07 W=1.19e-06 $X=2485 $Y=6020 $D=25
M9 Y 9 VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=3080 $Y=6020 $D=25
.ENDS
***************************************
.SUBCKT inv02 VSS VDD Y A
** N=4 EP=4 IP=0 FDC=2
M0 Y A VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1750 $D=19
M1 Y A VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=805 $Y=4970 $D=25
.ENDS
***************************************
.SUBCKT ALU_16Bit VSS VDD CB nBitOut[15] B[10] B[3] nBitOut[3] nBitOut[10] B[4] A[3] A[10] Control[1] nBitOut[9] A[9] Control[0] A[4] B[8] B[7] B[6] B[9]
+ nBitOut[7] nBitOut[4] nBitOut[6] B[11] A[7] A[6] B[0] B[13] B[5] A[0] A[8] nBitOut[5] nBitOut[11] A[11] nBitOut[8] A[5] A[12] A[13] nBitOut[12] nBitOut[13]
+ B[12] B[2] A[2] A[15] B[14] nBitOut[0] B[1] nBitOut[2] A[14] B[15] A[1] nBitOut[1] nBitOut[14]
** N=304 EP=53 IP=966 FDC=1138
M0 VSS B[0] 1 VSS nmos L=1.4e-07 W=3.5e-07 $X=46440 $Y=76000 $D=19
M1 3 B[0] VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=47035 $Y=75580 $D=19
M2 4 A[0] 3 VSS nmos L=1.4e-07 W=7.7e-07 $X=47455 $Y=75580 $D=19
M3 5 43 4 VSS nmos L=1.4e-07 W=7.7e-07 $X=48015 $Y=75580 $D=19
M4 VSS 1 5 VSS nmos L=1.4e-07 W=7.7e-07 $X=48435 $Y=75580 $D=19
M5 7 4 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=48995 $Y=75580 $D=19
M6 8 140 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=59940 $Y=47430 $D=19
M7 9 Control[1] 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=60360 $Y=47430 $D=19
M8 10 141 9 VSS nmos L=1.4e-07 W=1.19e-06 $X=60955 $Y=47010 $D=19
M9 11 Control[0] 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=61375 $Y=47010 $D=19
M10 VSS 202 11 VSS nmos L=1.4e-07 W=1.19e-06 $X=61795 $Y=47010 $D=19
M11 13 43 12 VSS nmos L=1.4e-07 W=7.7e-07 $X=62075 $Y=18860 $D=19
M12 VSS 207 13 VSS nmos L=1.4e-07 W=7.7e-07 $X=62495 $Y=18860 $D=19
M13 CB 207 14 VSS nmos L=1.4e-07 W=7.7e-07 $X=63615 $Y=18860 $D=19
M14 14 43 CB VSS nmos L=1.4e-07 W=7.7e-07 $X=64175 $Y=18860 $D=19
M15 VSS 12 14 VSS nmos L=1.4e-07 W=7.7e-07 $X=64735 $Y=18860 $D=19
M16 nBitOut[15] 211 16 VSS nmos L=1.4e-07 W=1.19e-06 $X=66485 $Y=47430 $D=19
M17 16 214 nBitOut[15] VSS nmos L=1.4e-07 W=1.19e-06 $X=67045 $Y=47430 $D=19
M18 16 19 18 VSS nmos L=1.4e-07 W=1.19e-06 $X=68165 $Y=47430 $D=19
M19 18 204 16 VSS nmos L=1.4e-07 W=1.19e-06 $X=68725 $Y=47430 $D=19
M20 VSS 219 18 VSS nmos L=1.4e-07 W=1.19e-06 $X=69285 $Y=47430 $D=19
M21 18 56 VSS VSS nmos L=1.4e-07 W=1.19e-06 $X=69845 $Y=47430 $D=19
M22 20 176 19 VSS nmos L=1.4e-07 W=9.1e-07 $X=72555 $Y=47010 $D=19
M23 VSS B[15] 20 VSS nmos L=1.4e-07 W=9.1e-07 $X=72975 $Y=47010 $D=19
M24 21 234 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=73570 $Y=47150 $D=19
M25 19 209 21 VSS nmos L=1.4e-07 W=7.7e-07 $X=73990 $Y=47150 $D=19
M26 VSS 66 19 VSS nmos L=1.4e-07 W=3.5e-07 $X=74585 $Y=47570 $D=19
M27 22 7 VSS VSS nmos L=1.4e-07 W=1.19e-06 $X=75905 $Y=75580 $D=19
M28 23 Control[1] 22 VSS nmos L=1.4e-07 W=1.19e-06 $X=76325 $Y=75580 $D=19
M29 24 229 23 VSS nmos L=1.4e-07 W=1.19e-06 $X=76745 $Y=75580 $D=19
M30 VDD B[0] 1 VDD pmos L=1.4e-07 W=7.7e-07 $X=46440 $Y=80060 $D=25
M31 25 B[0] VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=47035 $Y=80060 $D=25
M32 4 43 25 VDD pmos L=1.4e-07 W=1.54e-06 $X=47455 $Y=80060 $D=25
M33 26 A[0] 4 VDD pmos L=1.4e-07 W=1.54e-06 $X=48015 $Y=80060 $D=25
M34 VDD 1 26 VDD pmos L=1.4e-07 W=1.54e-06 $X=48435 $Y=80060 $D=25
M35 7 4 VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=48995 $Y=80060 $D=25
M36 9 140 27 VDD pmos L=1.4e-07 W=1.19e-06 $X=59555 $Y=51840 $D=25
M37 27 Control[1] 9 VDD pmos L=1.4e-07 W=1.19e-06 $X=60115 $Y=51840 $D=25
M38 VDD 141 27 VDD pmos L=1.4e-07 W=1.19e-06 $X=60675 $Y=51840 $D=25
M39 27 Control[0] VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=61235 $Y=51840 $D=25
M40 VDD 202 27 VDD pmos L=1.4e-07 W=1.19e-06 $X=61795 $Y=51840 $D=25
M41 12 43 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=62445 $Y=21835 $D=25
M42 VDD 207 12 VDD pmos L=1.4e-07 W=1.19e-06 $X=63005 $Y=21835 $D=25
M43 28 43 VDD VDD pmos L=1.4e-07 W=2.24e-06 $X=63635 $Y=21870 $D=25
M44 CB 207 28 VDD pmos L=1.4e-07 W=2.24e-06 $X=64125 $Y=21835 $D=25
M45 VDD 12 CB VDD pmos L=1.4e-07 W=1.19e-06 $X=64720 $Y=21870 $D=25
M46 29 211 VDD VDD pmos L=1.4e-07 W=2.52e-06 $X=67045 $Y=50510 $D=25
M47 nBitOut[15] 214 29 VDD pmos L=1.4e-07 W=2.52e-06 $X=67465 $Y=50510 $D=25
M48 30 19 nBitOut[15] VDD pmos L=1.4e-07 W=2.52e-06 $X=68025 $Y=50510 $D=25
M49 VDD 204 30 VDD pmos L=1.4e-07 W=2.52e-06 $X=68445 $Y=50510 $D=25
M50 31 219 VDD VDD pmos L=1.4e-07 W=2.52e-06 $X=69005 $Y=50510 $D=25
M51 nBitOut[15] 56 31 VDD pmos L=1.4e-07 W=2.52e-06 $X=69425 $Y=50510 $D=25
M52 VDD 176 32 VDD pmos L=1.4e-07 W=1.61e-06 $X=71785 $Y=51420 $D=25
M53 32 B[15] VDD VDD pmos L=1.4e-07 W=1.61e-06 $X=72345 $Y=51420 $D=25
M54 32 234 33 VDD pmos L=1.4e-07 W=1.61e-06 $X=73465 $Y=51420 $D=25
M55 33 209 32 VDD pmos L=1.4e-07 W=1.61e-06 $X=74025 $Y=51420 $D=25
M56 19 66 33 VDD pmos L=1.4e-07 W=1.61e-06 $X=74585 $Y=51420 $D=25
M57 VDD 7 24 VDD pmos L=1.4e-07 W=1.26e-06 $X=75765 $Y=80340 $D=25
M58 24 Control[1] VDD VDD pmos L=1.4e-07 W=1.26e-06 $X=76325 $Y=80340 $D=25
M59 VDD 229 24 VDD pmos L=1.4e-07 W=1.26e-06 $X=76885 $Y=80340 $D=25
X60 VSS VDD 37 B[10] inv01 $T=20 2965 0 0 $X=20 $Y=2965
X61 VSS VDD 41 36 inv01 $T=20 45820 0 0 $X=20 $Y=45820
X62 VSS VDD 38 B[3] inv01 $T=20 60105 0 0 $X=20 $Y=60105
X63 VSS VDD 67 49 inv01 $T=6390 88675 0 0 $X=6390 $Y=88675
X64 VSS VDD 54 59 inv01 $T=9330 60105 1 180 $X=7370 $Y=60105
X65 VSS VDD 42 71 inv01 $T=8350 31535 0 0 $X=8350 $Y=31535
X66 VSS VDD 53 68 inv01 $T=9330 2965 0 0 $X=9330 $Y=2965
X67 VSS VDD 74 61 inv01 $T=9330 45820 0 0 $X=9330 $Y=45820
X68 VSS VDD 73 B[4] inv01 $T=9330 60105 0 0 $X=9330 $Y=60105
X69 VSS VDD 99 B[6] inv01 $T=16680 88675 0 0 $X=16680 $Y=88675
X70 VSS VDD 88 B[9] inv01 $T=20110 17250 1 180 $X=18150 $Y=17250
X71 VSS VDD 106 B[7] inv01 $T=18150 31535 0 0 $X=18150 $Y=31535
X72 VSS VDD 110 102 inv01 $T=20110 17250 0 0 $X=20110 $Y=17250
X73 VSS VDD 117 83 inv01 $T=21580 45820 0 0 $X=21580 $Y=45820
X74 VSS VDD 114 121 inv01 $T=25500 31535 0 0 $X=25500 $Y=31535
X75 VSS VDD 105 120 inv01 $T=28930 88675 1 180 $X=26970 $Y=88675
X76 VSS VDD 129 B[13] inv01 $T=27460 17250 0 0 $X=27460 $Y=17250
X77 VSS VDD 130 B[8] inv01 $T=28440 60105 0 0 $X=28440 $Y=60105
X78 VSS VDD 133 B[11] inv01 $T=29910 2965 0 0 $X=29910 $Y=2965
X79 VSS VDD 76 136 inv01 $T=34320 31535 0 0 $X=34320 $Y=31535
X80 VSS VDD 115 96 inv01 $T=35300 60105 0 0 $X=35300 $Y=60105
X81 VSS VDD 150 122 inv01 $T=35790 17250 0 0 $X=35790 $Y=17250
X82 VSS VDD 148 138 inv01 $T=35790 74390 0 0 $X=35790 $Y=74390
X83 VSS VDD 66 56 inv01 $T=37260 60105 0 0 $X=37260 $Y=60105
X84 VSS VDD 151 157 inv01 $T=45590 74390 1 180 $X=43630 $Y=74390
X85 VSS VDD 132 75 inv01 $T=46080 45820 1 180 $X=44120 $Y=45820
X86 VSS VDD 178 169 inv01 $T=47060 60105 1 180 $X=45100 $Y=60105
X87 VSS VDD 177 163 inv01 $T=46080 45820 0 0 $X=46080 $Y=45820
X88 VSS VDD 46 72 inv01 $T=50000 74390 0 0 $X=50000 $Y=74390
X89 VSS VDD 153 B[5] inv01 $T=52940 31535 1 180 $X=50980 $Y=31535
X90 VSS VDD 181 B[12] inv01 $T=53920 17250 1 180 $X=51960 $Y=17250
X91 VSS VDD 172 187 inv01 $T=54900 31535 1 180 $X=52940 $Y=31535
X92 VSS VDD 149 164 inv01 $T=55880 17250 1 180 $X=53920 $Y=17250
X93 VSS VDD 190 139 inv01 $T=59800 88675 1 180 $X=57840 $Y=88675
X94 VSS VDD 200 B[2] inv01 $T=60780 60105 0 0 $X=60780 $Y=60105
X95 VSS VDD 204 A[15] inv01 $T=61760 31535 0 0 $X=61760 $Y=31535
X96 VSS VDD 179 182 inv01 $T=66170 17250 0 0 $X=66170 $Y=17250
X97 VSS VDD 216 B[1] inv01 $T=67150 88675 0 0 $X=67150 $Y=88675
X98 VSS VDD 221 193 inv01 $T=67640 74390 0 0 $X=67640 $Y=74390
X99 VSS VDD 220 B[14] inv01 $T=68130 2965 0 0 $X=68130 $Y=2965
X100 VSS VDD 219 B[15] inv01 $T=72050 31535 1 180 $X=70090 $Y=31535
X101 VSS VDD 202 7 inv01 $T=77930 60105 1 180 $X=75970 $Y=60105
X102 VSS VDD 231 209 inv01 $T=78910 31535 1 180 $X=76950 $Y=31535
X103 VSS VDD 208 233 inv01 $T=78910 31535 0 0 $X=78910 $Y=31535
X104 VSS VDD 199 226 inv01 $T=82975 74390 1 180 $X=81015 $Y=74390
X105 VSS VDD 239 217 inv01 $T=83810 17250 1 180 $X=81850 $Y=17250
X106 VSS VDD 141 A[0] 116 or02 $T=32850 74390 0 0 $X=32850 $Y=74390
X107 VSS VDD 238 7 229 or02 $T=81360 60105 0 0 $X=81360 $Y=60105
X108 VSS 64 VDD 71 41 nand02 $T=9330 45820 1 180 $X=6880 $Y=45820
X109 VSS 57 VDD 72 67 nand02 $T=10800 88675 1 180 $X=8350 $Y=88675
X110 VSS 81 VDD 59 74 nand02 $T=11290 60105 0 0 $X=11290 $Y=60105
X111 VSS 124 VDD 121 110 nand02 $T=25010 17250 0 0 $X=25010 $Y=17250
X112 VSS 125 VDD 120 117 nand02 $T=25990 60105 0 0 $X=25990 $Y=60105
X113 VSS 82 VDD 136 132 nand02 $T=32360 45820 1 180 $X=29910 $Y=45820
X114 VSS 158 VDD 68 150 nand02 $T=40200 17250 1 180 $X=37750 $Y=17250
X115 VSS 155 VDD 96 148 nand02 $T=37750 74390 0 0 $X=37750 $Y=74390
X116 VSS 183 VDD 164 177 nand02 $T=50490 45820 1 180 $X=48040 $Y=45820
X117 VSS 180 VDD 187 178 nand02 $T=52450 60105 1 180 $X=50000 $Y=60105
X118 VSS 185 VDD 157 190 nand02 $T=52450 88675 0 0 $X=52450 $Y=88675
X119 VSS 198 VDD Control[1] Control[0] nand02 $T=58820 2965 0 0 $X=58820 $Y=2965
X120 VSS 196 VDD 226 221 nand02 $T=72050 74390 1 180 $X=69600 $Y=74390
X121 VSS 214 VDD 207 Control[1] nand02 $T=72050 31535 0 0 $X=72050 $Y=31535
X122 VSS 218 VDD 233 231 nand02 $T=76950 31535 1 180 $X=74500 $Y=31535
X123 VSS 236 VDD 182 239 nand02 $T=79400 17250 0 0 $X=79400 $Y=17250
X124 VDD nBitOut[10] VSS 47 50 53 56 37 63 oai321 $T=1980 2965 0 0 $X=1980 $Y=2965
X125 VDD nBitOut[3] VSS 48 51 54 56 38 60 oai321 $T=1980 60105 0 0 $X=1980 $Y=60105
X126 VDD nBitOut[9] VSS 77 50 42 56 88 91 oai321 $T=12760 17250 0 0 $X=12760 $Y=17250
X127 VDD nBitOut[6] VSS 113 51 105 56 99 98 oai321 $T=24030 88675 1 180 $X=18640 $Y=88675
X128 VDD nBitOut[7] VSS 119 50 114 56 106 103 oai321 $T=25500 31535 1 180 $X=20110 $Y=31535
X129 VDD nBitOut[4] VSS 100 51 115 56 73 95 oai321 $T=25990 60105 1 180 $X=20600 $Y=60105
X130 VDD nBitOut[11] VSS 152 50 149 56 133 144 oai321 $T=40200 2965 1 180 $X=34810 $Y=2965
X131 VDD nBitOut[5] VSS 147 51 151 56 153 156 oai321 $T=35790 45820 0 0 $X=35790 $Y=45820
X132 VDD nBitOut[8] VSS 145 50 76 56 130 142 oai321 $T=39710 60105 0 0 $X=39710 $Y=60105
X133 VDD nBitOut[13] VSS 171 176 179 56 129 173 oai321 $T=51960 2965 1 180 $X=46570 $Y=2965
X134 VDD nBitOut[12] VSS 165 176 172 56 181 184 oai321 $T=46570 17250 0 0 $X=46570 $Y=17250
X135 VDD nBitOut[2] VSS 213 51 46 56 200 210 oai321 $T=65680 60105 0 0 $X=65680 $Y=60105
X136 VDD nBitOut[14] VSS 230 176 208 56 220 235 oai321 $T=82830 2965 1 180 $X=77440 $Y=2965
X137 VDD nBitOut[1] VSS 240 51 199 56 216 232 oai321 $T=84300 88675 1 180 $X=78910 $Y=88675
X138 VSS VDD 36 44 B[10] xor2 $T=20 31535 0 0 $X=20 $Y=31535
X139 VSS VDD 49 43 B[3] xor2 $T=20 74390 0 0 $X=20 $Y=74390
X140 VSS VDD 61 43 B[4] xor2 $T=1980 45820 0 0 $X=1980 $Y=45820
X141 VSS VDD 83 43 B[7] xor2 $T=18150 31535 1 180 $X=13250 $Y=31535
X142 VSS VDD 102 43 B[8] xor2 $T=16190 2965 0 0 $X=16190 $Y=2965
X143 VSS VDD 122 44 B[11] xor2 $T=21090 2965 0 0 $X=21090 $Y=2965
X144 VSS VDD 116 44 B[0] xor2 $T=27950 74390 1 180 $X=23050 $Y=74390
X145 VSS VDD 138 43 B[5] xor2 $T=27950 74390 0 0 $X=27950 $Y=74390
X146 VSS VDD 139 43 B[6] xor2 $T=28930 88675 0 0 $X=28930 $Y=88675
X147 VSS VDD 140 B[0] A[0] xor2 $T=30400 60105 0 0 $X=30400 $Y=60105
X148 VSS VDD 75 44 B[9] xor2 $T=36770 31535 0 0 $X=36770 $Y=31535
X149 VSS VDD 193 43 B[2] xor2 $T=52450 74390 0 0 $X=52450 $Y=74390
X150 VSS VDD 163 44 B[12] xor2 $T=58820 45820 1 180 $X=53920 $Y=45820
X151 VSS VDD 169 44 B[13] xor2 $T=67150 88675 1 180 $X=62250 $Y=88675
X152 VSS VDD 217 44 B[14] xor2 $T=63230 2965 0 0 $X=63230 $Y=2965
X153 VSS VDD 229 43 B[1] xor2 $T=71070 60105 0 0 $X=71070 $Y=60105
X154 VSS VDD 209 44 B[15] xor2 $T=83320 45820 1 180 $X=78420 $Y=45820
X155 47 VDD VSS 42 A[10] 36 nor03 $T=2960 17250 1 180 $X=20 $Y=17250
X156 48 VDD VSS 46 A[3] 49 nor03 $T=2960 88675 1 180 $X=20 $Y=88675
X157 77 VDD VSS 76 A[9] 75 nor03 $T=13250 31535 1 180 $X=10310 $Y=31535
X158 100 VDD VSS 54 A[4] 61 nor03 $T=17660 60105 0 0 $X=17660 $Y=60105
X159 119 VDD VSS 105 A[7] 83 nor03 $T=26480 45820 1 180 $X=23540 $Y=45820
X160 145 VDD VSS 114 A[8] 102 nor03 $T=32850 17250 0 0 $X=32850 $Y=17250
X161 152 VDD VSS 53 A[11] 122 nor03 $T=43140 2965 1 180 $X=40200 $Y=2965
X162 113 VDD VSS 151 A[6] 139 nor03 $T=44120 88675 1 180 $X=41180 $Y=88675
X163 165 VDD VSS 149 A[12] 163 nor03 $T=44610 31535 1 180 $X=41670 $Y=31535
X164 171 VDD VSS 172 A[13] 169 nor03 $T=46570 17250 1 180 $X=43630 $Y=17250
X165 147 VDD VSS 115 A[5] 138 nor03 $T=47060 60105 0 0 $X=47060 $Y=60105
X166 211 VDD VSS 208 A[15] 209 nor03 $T=63720 31535 0 0 $X=63720 $Y=31535
X167 213 VDD VSS 199 A[2] 193 nor03 $T=64700 74390 0 0 $X=64700 $Y=74390
X168 230 VDD VSS 179 A[14] 217 nor03 $T=70090 2965 0 0 $X=70090 $Y=2965
X169 240 VDD VSS 7 A[1] 229 nor03 $T=77930 74390 0 0 $X=77930 $Y=74390
X170 VSS VDD 59 49 46 A[3] 57 aoi22 $T=2960 88675 0 0 $X=2960 $Y=88675
X171 VSS VDD 68 36 42 A[10] 64 aoi22 $T=4920 31535 0 0 $X=4920 $Y=31535
X172 VSS VDD 71 75 76 A[9] 82 aoi22 $T=11290 45820 0 0 $X=11290 $Y=45820
X173 VSS VDD 96 61 54 A[4] 81 aoi22 $T=14230 60105 0 0 $X=14230 $Y=60105
X174 VSS VDD 121 83 105 A[7] 125 aoi22 $T=26480 45820 0 0 $X=26480 $Y=45820
X175 VSS VDD 136 102 114 A[8] 124 aoi22 $T=29420 17250 0 0 $X=29420 $Y=17250
X176 VSS VDD 164 122 53 A[11] 158 aoi22 $T=40200 17250 0 0 $X=40200 $Y=17250
X177 VSS VDD 157 138 115 A[5] 155 aoi22 $T=43630 74390 1 180 $X=40200 $Y=74390
X178 VSS VDD 182 169 172 A[13] 180 aoi22 $T=47550 31535 0 0 $X=47550 $Y=31535
X179 VSS VDD 120 139 151 A[6] 185 aoi22 $T=49020 88675 0 0 $X=49020 $Y=88675
X180 VSS VDD 187 163 149 A[12] 183 aoi22 $T=50490 45820 0 0 $X=50490 $Y=45820
X181 VSS VDD 72 193 199 A[2] 196 aoi22 $T=60780 74390 1 180 $X=57350 $Y=74390
X182 VSS VDD 207 209 208 A[15] 218 aoi22 $T=66660 31535 0 0 $X=66660 $Y=31535
X183 VSS VDD 233 217 179 A[14] 236 aoi22 $T=75970 17250 0 0 $X=75970 $Y=17250
X184 VSS VDD 226 229 7 A[1] 238 aoi22 $T=77930 60105 0 0 $X=77930 $Y=60105
X185 VSS VDD 58 Control[1] 71 nor02ii $T=12760 17250 1 180 $X=9820 $Y=17250
X186 VSS VDD 65 Control[1] 72 nor02ii $T=13740 88675 1 180 $X=10800 $Y=88675
X187 VSS VDD 78 Control[0] Control[1] nor02ii $T=16190 2965 1 180 $X=13250 $Y=2965
X188 VSS VDD 85 Control[1] 59 nor02ii $T=13740 88675 0 0 $X=13740 $Y=88675
X189 VSS VDD 92 Control[1] 120 nor02ii $T=26970 88675 1 180 $X=24030 $Y=88675
X190 VSS VDD 127 Control[1] 121 nor02ii $T=30400 31535 1 180 $X=27460 $Y=31535
X191 VSS VDD 137 Control[1] 136 nor02ii $T=35300 45820 1 180 $X=32360 $Y=45820
X192 VSS VDD 143 Control[1] 157 nor02ii $T=40690 88675 1 180 $X=37750 $Y=88675
X193 VSS VDD 175 Control[1] 68 nor02ii $T=43140 2965 0 0 $X=43140 $Y=2965
X194 VSS VDD 191 Control[1] 96 nor02ii $T=52450 60105 0 0 $X=52450 $Y=60105
X195 VSS VDD 170 Control[1] 187 nor02ii $T=57840 88675 1 180 $X=54900 $Y=88675
X196 VSS VDD 194 Control[1] 164 nor02ii $T=61760 31535 1 180 $X=58820 $Y=31535
X197 VSS VDD 223 Control[1] 182 nor02ii $T=68130 17250 0 0 $X=68130 $Y=17250
X198 VSS VDD 203 Control[1] 226 nor02ii $T=74990 74390 1 180 $X=72050 $Y=74390
X199 VSS VDD 234 Control[1] 233 nor02ii $T=75480 45820 0 0 $X=75480 $Y=45820
X200 VSS 63 VDD A[10] 66 62 oai21 $T=6880 17250 0 0 $X=6880 $Y=17250
X201 VSS 60 VDD A[3] 66 70 oai21 $T=11780 74390 1 180 $X=8840 $Y=74390
X202 VSS 95 VDD A[4] 66 89 oai21 $T=19620 74390 1 180 $X=16680 $Y=74390
X203 VSS 103 VDD A[7] 66 84 oai21 $T=21580 45820 1 180 $X=18640 $Y=45820
X204 VSS 98 VDD A[6] 66 112 oai21 $T=23050 74390 1 180 $X=20110 $Y=74390
X205 VSS 91 VDD A[9] 66 118 oai21 $T=22070 17250 0 0 $X=22070 $Y=17250
X206 VSS 142 VDD A[8] 66 131 oai21 $T=31870 2965 0 0 $X=31870 $Y=2965
X207 VSS 156 VDD A[5] 66 161 oai21 $T=44120 45820 1 180 $X=41180 $Y=45820
X208 VSS 173 VDD A[13] 66 167 oai21 $T=44610 31535 0 0 $X=44610 $Y=31535
X209 VSS 144 VDD A[11] 66 192 oai21 $T=55880 2965 0 0 $X=55880 $Y=2965
X210 VSS 184 VDD A[12] 66 195 oai21 $T=56370 17250 0 0 $X=56370 $Y=17250
X211 VSS nBitOut[0] VDD 9 202 Control[1] oai21 $T=62740 45820 0 0 $X=62740 $Y=45820
X212 VSS 210 VDD A[2] 66 206 oai21 $T=65680 60105 1 180 $X=62740 $Y=60105
X213 VSS 227 VDD 24 216 Control[1] oai21 $T=74010 88675 1 180 $X=71070 $Y=88675
X214 VSS 232 VDD A[1] 66 227 oai21 $T=76950 88675 1 180 $X=74010 $Y=88675
X215 VSS 235 VDD A[14] 66 228 oai21 $T=74500 2965 0 0 $X=74500 $Y=2965
X216 VSS VDD 62 B[10] 36 58 50 ao22 $T=2960 17250 0 0 $X=2960 $Y=17250
X217 VSS VDD 70 B[3] 49 65 51 ao22 $T=4920 74390 0 0 $X=4920 $Y=74390
X218 VSS VDD 89 B[4] 61 85 51 ao22 $T=12760 74390 0 0 $X=12760 $Y=74390
X219 VSS VDD 84 B[7] 83 92 50 ao22 $T=18640 45820 1 180 $X=14720 $Y=45820
X220 VSS VDD 131 B[8] 102 127 50 ao22 $T=25990 2965 0 0 $X=25990 $Y=2965
X221 VSS VDD 118 B[9] 75 137 50 ao22 $T=34320 31535 1 180 $X=30400 $Y=31535
X222 VSS VDD 112 B[6] 139 143 50 ao22 $T=37750 88675 1 180 $X=33830 $Y=88675
X223 VSS VDD 167 B[13] 169 170 176 ao22 $T=48040 88675 1 180 $X=44120 $Y=88675
X224 VSS VDD 192 B[11] 122 175 176 ao22 $T=51960 2965 0 0 $X=51960 $Y=2965
X225 VSS VDD 195 B[12] 163 194 176 ao22 $T=54900 31535 0 0 $X=54900 $Y=31535
X226 VSS VDD 161 B[5] 138 191 51 ao22 $T=56860 60105 0 0 $X=56860 $Y=60105
X227 VSS VDD 206 B[2] 193 203 51 ao22 $T=60780 74390 0 0 $X=60780 $Y=74390
X228 VSS VDD 228 B[14] 217 223 176 ao22 $T=72050 17250 0 0 $X=72050 $Y=17250
X229 VSS VDD 50 Control[1] inv02 $T=9330 2965 1 180 $X=7370 $Y=2965
X230 VSS VDD 56 78 inv02 $T=13250 2965 1 180 $X=11290 $Y=2965
X231 VSS VDD 44 198 inv02 $T=59310 17250 0 0 $X=59310 $Y=17250
X232 VSS VDD 51 Control[1] inv02 $T=59800 88675 0 0 $X=59800 $Y=88675
X233 VSS VDD 43 198 inv02 $T=63230 2965 1 180 $X=61270 $Y=2965
X234 VSS VDD 176 Control[1] inv02 $T=69110 88675 0 0 $X=69110 $Y=88675
.ENDS
***************************************
