* Example circuit file for simulating PEX

.OPTION DOTNODE
.HIER /

.INCLUDE "/home/bxk5113/Pyxis_SPT_HEP/ic_projects/Pyxis_SPT/digicdesign/ALU_16Bit/ALU_16Bit.cal/ALU_16Bit.pex.netlist"

.LIB /home/bxk5113/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT

* - Instantiate your parasitic netlist and add the load capacitor
** FORMAT :
* XLAYOUT [all inputs as listed by the ".subckt" line in the included netlist, in the order that they appear there] [name of the subcircuit as listed in the included netlist]
XLAYOUT CB NBITOUT[15] NBITOUT[14] NBITOUT[13] NBITOUT[12] NBITOUT[11] NBITOUT[10] NBITOUT[9] NBITOUT[8] NBITOUT[7] NBITOUT[6] NBITOUT[5] NBITOUT[4] NBITOUT[3] NBITOUT[2] NBITOUT[1] NBITOUT[0] A[15] A[14] A[13] A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[15] B[14] B[13] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CONTROL[1] CONTROL[0] ALU_16Bit

* Output Capactitance
C_CB CB 0 120f
C_NBITOUT[15] NBITOUT[15] 0 120f
C_NBITOUT[14] NBITOUT[14] 0 120f
C_NBITOUT[13] NBITOUT[13] 0 120f
C_NBITOUT[12] NBITOUT[12] 0 120f
C_NBITOUT[11] NBITOUT[11] 0 120f
C_NBITOUT[10] NBITOUT[10] 0 120f
C_NBITOUT[9] NBITOUT[9] 0 120f
C_NBITOUT[8] NBITOUT[8] 0 120f
C_NBITOUT[7] NBITOUT[7] 0 120f
C_NBITOUT[6] NBITOUT[6] 0 120f
C_NBITOUT[5] NBITOUT[5] 0 120f
C_NBITOUT[4] NBITOUT[4] 0 120f
C_NBITOUT[3] NBITOUT[3] 0 120f
C_NBITOUT[2] NBITOUT[2] 0 120f
C_NBITOUT[1] NBITOUT[1] 0 120f
C_NBITOUT[0] NBITOUT[0] 0 120f


* - Analysis Setup - DC sweep
* FORMAT : .DC [name] [low] [high] [step]
*.DC VFORCE__A 0 1.2 0.01

* - Analysis Setup - Trans
* FORMAT : .TRAN [start time] [end time] [time step]
.TRAN 0 400n 0.001n

* --- Forces
* FORMAT -- PULSE : [name] [port] [reference (0 means ground)] PULSE [low] [high] [delay] [fall time] [rise time] [pulse width] [period]
*
* FORMAT -- DC    : [name] [port] [reference (0 means ground)] DC [voltage]
*

VFORCE__C1 CONTROL[1] 0 PULSE (0 1.08 40n 0.1n 0.1n 40n 80n)
VFORCE__C0 CONTROL[0] 0 PULSE (0 1.08 20n 0.1n 0.1n 20n 40n)

VFORCE__VDD VDD 0 DC 1.08
VFORCE__VSS VSS 0 DC 0

VFORCE__A[0] A[0] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[1] A[1] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011000 R
VFORCE__A[2] A[2] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[3] A[3] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011000 R
VFORCE__A[4] A[4] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[5] A[5] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011000 R
VFORCE__A[6] A[6] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[7] A[7] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[8] A[8] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[9] A[9] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[10] A[10] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011000 R
VFORCE__A[11] A[11] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011000 R
VFORCE__A[12] A[12] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[13] A[13] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011001 R
VFORCE__A[14] A[14] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011000 R
VFORCE__A[15] A[15] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011101 R
VFORCE__B[0] B[0] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[1] B[1] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010100 R
VFORCE__B[2] B[2] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010100 R
VFORCE__B[3] B[3] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010100 R
VFORCE__B[4] B[4] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[5] B[5] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010100 R
VFORCE__B[6] B[6] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010100 R
VFORCE__B[7] B[7] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[8] B[8] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[9] B[9] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[10] B[10] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[11] B[11] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010100 R
VFORCE__B[12] B[12] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[13] B[13] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[14] B[14] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 010101 R
VFORCE__B[15] B[15] 0 PBIT 0 1.08 0 0 0.01n 0 0.01n 80n 011111 R





* --- Waveform Outputs
.PLOT TRAN V(CB)
.PLOT TRAN V(NBITOUT[15])
.PLOT TRAN V(NBITOUT[14])
.PLOT TRAN V(NBITOUT[13])
.PLOT TRAN V(NBITOUT[12])
.PLOT TRAN V(NBITOUT[11])
.PLOT TRAN V(NBITOUT[10])
.PLOT TRAN V(NBITOUT[9])
.PLOT TRAN V(NBITOUT[8])
.PLOT TRAN V(NBITOUT[7])
.PLOT TRAN V(NBITOUT[6])
.PLOT TRAN V(NBITOUT[5])
.PLOT TRAN V(NBITOUT[4])
.PLOT TRAN V(NBITOUT[3])
.PLOT TRAN V(NBITOUT[2])
.PLOT TRAN V(NBITOUT[1])
.PLOT TRAN V(NBITOUT[0])
.PLOT TRAN V(A[15])
.PLOT TRAN V(A[14])
.PLOT TRAN V(A[13])
.PLOT TRAN V(A[12])
.PLOT TRAN V(A[11])
.PLOT TRAN V(A[10])
.PLOT TRAN V(A[9])
.PLOT TRAN V(A[8])
.PLOT TRAN V(A[7])
.PLOT TRAN V(A[6])
.PLOT TRAN V(A[5])
.PLOT TRAN V(A[4])
.PLOT TRAN V(A[3])
.PLOT TRAN V(A[2])
.PLOT TRAN V(A[1])
.PLOT TRAN V(A[0])
.PLOT TRAN V(B[15])
.PLOT TRAN V(B[14])
.PLOT TRAN V(B[13])
.PLOT TRAN V(B[12])
.PLOT TRAN V(B[11])
.PLOT TRAN V(B[10])
.PLOT TRAN V(B[9])
.PLOT TRAN V(B[8])
.PLOT TRAN V(B[7])
.PLOT TRAN V(B[6])
.PLOT TRAN V(B[5])
.PLOT TRAN V(B[4])
.PLOT TRAN V(B[3])
.PLOT TRAN V(B[2])
.PLOT TRAN V(B[1])
.PLOT TRAN V(B[0])
.PLOT TRAN V(CONTROL[1])
.PLOT TRAN V(CONTROL[0])


* --- Params
.TEMP 125

* --- Power Measurement
.measure tran static_pwr AVG power from=90ns to=150ns
.measure tran inst_pwr MAX power from=90ns to=150ns

