* SPICE NETLIST
***************************************

.SUBCKT mimcap_g13 plus minus
.ENDS
***************************************
.SUBCKT spiral_inductor_lvs pos neg
.ENDS
***************************************
.SUBCKT mirroradder GROUND VDD Cout NS S B A Cin
** N=19 EP=8 IP=0 FDC=28
* PORT GROUND GROUND 4485 -1300 metal1
* PORT VDD VDD 4485 10010 metal1
* PORT Cout Cout 2730 3900 metal2
* PORT NS NS 7410 910 metal1
* PORT S S 10790 780 metal1
* PORT B B -1560 2470 metal2
* PORT A A -390 1820 metal2
* PORT Cin Cin 780 3380 metal2
M0 GROUND B 1 GROUND nmos L=1.3e-07 W=5.2e-07 $X=-1560 $Y=1040 $D=19
M1 3 B GROUND GROUND nmos L=1.3e-07 W=5.2e-07 $X=-650 $Y=1040 $D=19
M2 4 A 3 GROUND nmos L=1.3e-07 W=5.2e-07 $X=-130 $Y=1040 $D=19
M3 1 Cin 4 GROUND nmos L=1.3e-07 W=5.2e-07 $X=780 $Y=1040 $D=19
M4 GROUND A 1 GROUND nmos L=1.3e-07 W=5.2e-07 $X=1430 $Y=1040 $D=19
M5 Cout 4 GROUND GROUND nmos L=1.3e-07 W=2.6e-07 $X=2340 $Y=1170 $D=19
M6 7 Cin GROUND GROUND nmos L=1.3e-07 W=5.2e-07 $X=4160 $Y=1040 $D=19
M7 GROUND B 7 GROUND nmos L=1.3e-07 W=5.2e-07 $X=5070 $Y=1040 $D=19
M8 7 A GROUND GROUND nmos L=1.3e-07 W=5.2e-07 $X=5980 $Y=1040 $D=19
M9 NS 4 7 GROUND nmos L=1.3e-07 W=5.2e-07 $X=7020 $Y=1040 $D=19
M10 9 Cin NS GROUND nmos L=1.3e-07 W=7.8e-07 $X=7930 $Y=780 $D=19
M11 10 B 9 GROUND nmos L=1.3e-07 W=7.8e-07 $X=8840 $Y=780 $D=19
M12 GROUND A 10 GROUND nmos L=1.3e-07 W=7.8e-07 $X=9490 $Y=780 $D=19
M13 S NS GROUND GROUND nmos L=1.3e-07 W=2.6e-07 $X=10400 $Y=1170 $D=19
M14 VDD B 12 VDD pmos L=1.3e-07 W=1.04e-06 $X=-1560 $Y=6370 $D=25
M15 13 B VDD VDD pmos L=1.3e-07 W=1.04e-06 $X=-650 $Y=6370 $D=25
M16 4 A 13 VDD pmos L=1.3e-07 W=1.04e-06 $X=-130 $Y=6370 $D=25
M17 12 Cin 4 VDD pmos L=1.3e-07 W=1.04e-06 $X=780 $Y=6370 $D=25
M18 VDD A 12 VDD pmos L=1.3e-07 W=1.04e-06 $X=1430 $Y=6370 $D=25
M19 Cout 4 VDD VDD pmos L=1.3e-07 W=5.2e-07 $X=2340 $Y=6630 $D=25
M20 14 Cin VDD VDD pmos L=1.3e-07 W=1.04e-06 $X=4160 $Y=6370 $D=25
M21 VDD B 14 VDD pmos L=1.3e-07 W=1.04e-06 $X=5070 $Y=6370 $D=25
M22 14 A VDD VDD pmos L=1.3e-07 W=1.04e-06 $X=5980 $Y=6370 $D=25
M23 NS 4 14 VDD pmos L=1.3e-07 W=1.04e-06 $X=7020 $Y=6370 $D=25
M24 15 Cin NS VDD pmos L=1.3e-07 W=1.56e-06 $X=7930 $Y=6370 $D=25
M25 16 B 15 VDD pmos L=1.3e-07 W=1.56e-06 $X=8840 $Y=6370 $D=25
M26 VDD A 16 VDD pmos L=1.3e-07 W=1.56e-06 $X=9490 $Y=6370 $D=25
M27 S NS VDD VDD pmos L=1.3e-07 W=5.2e-07 $X=10400 $Y=6630 $D=25
.ENDS
***************************************
