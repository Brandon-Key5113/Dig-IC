//
// Verilog description for cell MAC, 
// Fri Nov 22 17:41:19 2019
//
// LeonardoSpectrum Level 3, 2008b.3 
//


module MAC ( A, B, clk, WE, reset, RegOut ) ;

    input [15:0]A ;
    input [15:0]B ;
    input clk ;
    input WE ;
    input reset ;
    output [31:0]RegOut ;

    wire MultA_15, MultA_14, MultA_13, MultA_12, MultA_11, MultA_10, MultA_9, 
         MultA_8, MultA_7, MultA_6, MultA_5, MultA_4, MultA_3, MultA_2, MultA_1, 
         MultA_0, MultB_15, MultB_14, MultB_13, MultB_12, MultB_11, MultB_10, 
         MultB_9, MultB_8, MultB_7, MultB_6, MultB_5, MultB_4, MultB_3, MultB_2, 
         MultB_1, MultB_0, Product_31, Product_30, Product_29, Product_28, 
         Product_27, Product_26, Product_25, Product_24, Product_23, Product_22, 
         Product_21, Product_20, Product_19, Product_18, Product_17, Product_16, 
         Product_0, adderB_31, adderB_30, adderB_29, adderB_28, adderB_27, 
         adderB_26, adderB_25, adderB_24, adderB_23, adderB_22, adderB_21, 
         adderB_20, adderB_19, adderB_18, adderB_17, adderB_16, adderB_15, 
         adderB_14, adderB_13, adderB_12, adderB_11, adderB_10, adderB_9, 
         adderB_8, adderB_7, adderB_6, adderB_5, adderB_4, adderB_3, adderB_2, 
         adderB_1, adderB_0, adderOut_31, adderOut_30, adderOut_29, adderOut_28, 
         adderOut_27, adderOut_26, adderOut_25, adderOut_24, adderOut_23, 
         adderOut_22, adderOut_21, adderOut_20, adderOut_19, adderOut_18, 
         adderOut_17, adderOut_16, adderOut_15, adderOut_14, adderOut_13, 
         adderOut_12, adderOut_11, adderOut_10, adderOut_9, adderOut_8, 
         adderOut_7, adderOut_6, adderOut_5, adderOut_4, adderOut_3, adderOut_2, 
         adderOut_1, adderOut_0, ADD1_c_array_30, ADD1_c_array_29, 
         ADD1_c_array_28, ADD1_c_array_27, ADD1_c_array_26, ADD1_c_array_25, 
         ADD1_c_array_24, ADD1_c_array_23, ADD1_c_array_22, ADD1_c_array_21, 
         ADD1_c_array_20, ADD1_c_array_19, ADD1_c_array_18, ADD1_c_array_17, 
         ADD1_c_array_16, ADD1_c_array_15, ADD1_c_array_14, ADD1_c_array_13, 
         ADD1_c_array_12, ADD1_c_array_11, ADD1_c_array_10, ADD1_c_array_9, 
         ADD1_c_array_8, ADD1_c_array_7, ADD1_c_array_6, ADD1_c_array_5, 
         ADD1_c_array_4, ADD1_c_array_3, ADD1_c_array_2, ADD1_c_array_1, 
         ADD1_c_array_0, Product_1, Product_2, Product_3, Product_4, Product_5, 
         Product_6, Product_7, Product_8, Product_9, Product_10, Product_11, 
         Product_12, Product_13, Product_14, Product_15, MULT1_F_1024, PWR, nx14, 
         nx22, nx30, nx32, nx38, nx46, nx54, nx62, nx64, nx66, nx68, nx74, nx82, 
         nx90, nx98, nx106, nx108, nx110, nx112, nx114, nx116, nx122, nx130, 
         nx138, nx146, nx154, nx162, nx164, nx166, nx168, nx170, nx172, nx174, 
         nx176, nx182, nx190, nx198, nx206, nx214, nx222, nx230, nx232, nx234, 
         nx236, nx238, nx240, nx242, nx244, nx246, nx248, nx254, nx262, nx270, 
         nx278, nx286, nx294, nx302, nx310, nx312, nx314, nx316, nx318, nx320, 
         nx322, nx324, nx326, nx328, nx330, nx332, nx338, nx346, nx354, nx362, 
         nx370, nx378, nx386, nx394, nx402, nx404, nx406, nx408, nx410, nx412, 
         nx414, nx416, nx418, nx420, nx422, nx424, nx426, nx428, nx434, nx442, 
         nx450, nx458, nx466, nx474, nx482, nx490, nx498, nx506, nx508, nx510, 
         nx512, nx514, nx516, nx518, nx520, nx522, nx524, nx526, nx528, nx530, 
         nx532, nx534, nx536, nx542, nx550, nx558, nx566, nx574, nx582, nx590, 
         nx598, nx606, nx614, nx622, nx624, nx626, nx628, nx630, nx632, nx634, 
         nx636, nx638, nx640, nx642, nx644, nx646, nx648, nx650, nx652, nx654, 
         nx656, nx662, nx670, nx678, nx686, nx694, nx702, nx710, nx718, nx726, 
         nx734, nx742, nx750, nx752, nx754, nx756, nx758, nx760, nx762, nx764, 
         nx766, nx768, nx770, nx772, nx774, nx776, nx778, nx780, nx782, nx784, 
         nx786, nx788, nx794, nx802, nx810, nx818, nx826, nx834, nx842, nx850, 
         nx858, nx866, nx874, nx882, nx890, nx892, nx894, nx896, nx898, nx900, 
         nx902, nx904, nx906, nx908, nx910, nx912, nx914, nx916, nx918, nx920, 
         nx922, nx924, nx926, nx928, nx930, nx932, nx938, nx946, nx954, nx962, 
         nx970, nx978, nx986, nx994, nx1002, nx1010, nx1018, nx1026, nx1034, 
         nx1042, nx1044, nx1046, nx1048, nx1050, nx1052, nx1054, nx1056, nx1058, 
         nx1060, nx1062, nx1064, nx1066, nx1068, nx1070, nx1072, nx1074, nx1076, 
         nx1078, nx1080, nx1082, nx1084, nx1086, nx1088, nx1094, nx1102, nx1110, 
         nx1118, nx1126, nx1134, nx1142, nx1150, nx1158, nx1166, nx1174, nx1182, 
         nx1190, nx1198, nx1206, nx1208, nx1210, nx1212, nx1214, nx1216, nx1218, 
         nx1220, nx1222, nx1224, nx1226, nx1228, nx1230, nx1232, nx1234, nx1236, 
         nx1238, nx1240, nx1242, nx1244, nx1246, nx1248, nx1250, nx1252, nx1254, 
         nx1256, nx1262, nx1374, nx1376, nx1446, nx1454, nx1462, nx1470, nx1478, 
         nx1486, nx1494, nx1502, nx1510, nx1518, nx1526, nx1534, nx1542, nx1550, 
         nx1556, nx1558, nx1564, nx1566, nx1572, nx1574, nx1580, nx1582, nx1588, 
         nx1590, nx1596, nx1598, nx1604, nx1606, nx1612, nx1620, nx1636, nx1644, 
         nx1652, nx1668, nx1676, nx1684, nx1700, nx1708, nx1716, nx1718, nx1720, 
         nx1722, nx1732, nx1734, nx1736, nx1738, nx1748, nx1750, nx1752, nx1754, 
         nx1764, nx1766, nx1780, nx1788, nx1812, nx1820, nx1844, nx1852, nx1876, 
         nx1878, nx1892, nx1894, nx1908, nx1910, nx1920, nx1936, nx1944, nx1952, 
         nx1960, nx1968, nx1976, nx1984, nx2000, nx2008, nx2010, nx2020, nx2022, 
         nx2028, nx2030, nx2032, nx2034, nx2040, nx2042, nx2056, nx2064, nx2080, 
         nx2088, nx2096, nx2104, nx2120, nx2128, nx2140, nx2142, nx2152, nx2154, 
         nx2156, nx2158, nx2160, nx2162, nx2172, nx2174, nx2180, nx2188, nx2196, 
         nx2204, nx2212, nx2220, nx2228, nx2236, nx2244, nx2252, nx2254, nx2256, 
         nx2258, nx2264, nx2266, nx2268, nx2270, nx2272, nx2274, nx2276, nx2278, 
         nx2284, nx2286, nx2300, nx2308, nx2316, nx2324, nx2332, nx2340, nx2364, 
         nx2366, nx2368, nx2370, nx2372, nx2374, nx2376, nx2378, nx2380, nx2382, 
         nx2392, nx2440, nx2448, nx2450, nx2480, nx2488, nx2496, nx2504, nx2512, 
         nx2520, nx2532, nx2534, nx2540, nx2542, nx2548, nx2550, nx2556, nx2564, 
         nx2580, nx2588, nx2596, nx2598, nx2600, nx2602, nx2612, nx2614, nx2628, 
         nx2636, nx2660, nx2662, nx2672, nx2688, nx2696, nx2698, nx2712, nx2720, 
         nx2732, nx2734, nx2740, nx2748, nx2750, nx2788, nx2796, nx2804, nx2812, 
         nx2820, nx2828, nx2836, nx2844, nx2852, nx2860, nx497, nx501, nx505, 
         nx509, nx513, nx517, nx521, nx525, nx529, nx533, nx537, nx541, nx545, 
         nx549, nx553, nx557, nx559, nx565, nx567, nx569, nx571, nx575, nx581, 
         nx583, nx585, nx587, nx589, nx593, nx597, nx601, nx607, nx609, nx611, 
         nx619, nx621, nx623, nx625, nx629, nx633, nx637, nx641, nx647, nx653, 
         nx655, nx661, nx663, nx665, nx667, nx671, nx675, nx679, nx683, nx689, 
         nx693, nx699, nx705, nx707, nx713, nx715, nx717, nx719, nx723, nx727, 
         nx731, nx735, nx741, nx745, nx751, nx755, nx761, nx767, nx769, nx775, 
         nx777, nx779, nx781, nx785, nx789, nx793, nx797, nx803, nx807, nx813, 
         nx817, nx823, nx827, nx833, nx839, nx841, nx847, nx849, nx851, nx853, 
         nx857, nx861, nx865, nx869, nx875, nx879, nx885, nx889, nx895, nx899, 
         nx905, nx909, nx915, nx921, nx923, nx929, nx931, nx933, nx935, nx939, 
         nx943, nx947, nx951, nx957, nx961, nx967, nx971, nx977, nx981, nx987, 
         nx991, nx997, nx1001, nx1007, nx1013, nx1015, nx1021, nx1023, nx1025, 
         nx1027, nx1031, nx1035, nx1039, nx1043, nx1049, nx1053, nx1059, nx1063, 
         nx1069, nx1073, nx1079, nx1083, nx1089, nx1093, nx1099, nx1103, nx1109, 
         nx1115, nx1117, nx1123, nx1125, nx1127, nx1129, nx1133, nx1137, nx1141, 
         nx1145, nx1151, nx1155, nx1161, nx1165, nx1171, nx1175, nx1181, nx1185, 
         nx1191, nx1195, nx1201, nx1205, nx1211, nx1215, nx1221, nx1227, nx1229, 
         nx1235, nx1237, nx1239, nx1241, nx1245, nx1249, nx1253, nx1257, nx1263, 
         nx1267, nx1273, nx1277, nx1283, nx1287, nx1293, nx1297, nx1303, nx1307, 
         nx1313, nx1317, nx1323, nx1327, nx1333, nx1337, nx1343, nx1349, nx1351, 
         nx1357, nx1359, nx1361, nx1363, nx1367, nx1371, nx1375, nx1379, nx1385, 
         nx1389, nx1395, nx1399, nx1405, nx1409, nx1415, nx1419, nx1425, nx1429, 
         nx1435, nx1439, nx1445, nx1449, nx1455, nx1459, nx1465, nx1469, nx1475, 
         nx1481, nx1483, nx1489, nx1491, nx1493, nx1495, nx1499, nx1503, nx1507, 
         nx1511, nx1517, nx1521, nx1527, nx1531, nx1537, nx1541, nx1547, nx1551, 
         nx1557, nx1561, nx1567, nx1571, nx1577, nx1581, nx1587, nx1591, nx1597, 
         nx1601, nx1607, nx1611, nx1617, nx1623, nx1625, nx1631, nx1633, nx1635, 
         nx1639, nx1645, nx1651, nx1657, nx1663, nx1669, nx1675, nx1681, nx1687, 
         nx1693, nx1697, nx1701, nx1705, nx1709, nx1715, nx1717, nx1719, nx1721, 
         nx1723, nx1725, nx1727, nx1729, nx1733, nx1735, nx1737, nx1739, nx1743, 
         nx1745, nx1747, nx1749, nx1753, nx1755, nx1757, nx1759, nx1763, nx1765, 
         nx1767, nx1769, nx1773, nx1775, nx1777, nx1779, nx1783, nx1785, nx1787, 
         nx1789, nx1793, nx1795, nx1797, nx1799, nx1803, nx1805, nx1807, nx1809, 
         nx1813, nx1815, nx1817, nx1819, nx1823, nx1825, nx1827, nx1829, nx1833, 
         nx1835, nx1837, nx1839, nx1843, nx1845, nx1847, nx1849, nx1853, nx1857, 
         nx1859, nx1873, nx1879, nx1881, nx1883, nx1889, nx1895, nx1897, nx1899, 
         nx1905, nx1911, nx1913, nx1915, nx1921, nx1927, nx1929, nx1931, nx1937, 
         nx1943, nx1945, nx1947, nx1953, nx1959, nx1961, nx1963, nx1969, nx1975, 
         nx1977, nx1979, nx1983, nx1987, nx1993, nx1995, nx1997, nx1999, nx2001, 
         nx2003, nx2005, nx2007, nx2011, nx2015, nx2019, nx2023, nx2029, nx2031, 
         nx2033, nx2035, nx2037, nx2039, nx2041, nx2043, nx2047, nx2051, nx2055, 
         nx2059, nx2065, nx2067, nx2069, nx2071, nx2073, nx2075, nx2077, nx2079, 
         nx2083, nx2087, nx2091, nx2095, nx2099, nx2103, nx2107, nx2109, nx2111, 
         nx2115, nx2123, nx2129, nx2131, nx2133, nx2135, nx2137, nx2139, nx2141, 
         nx2143, nx2147, nx2149, nx2151, nx2155, nx2163, nx2169, nx2171, nx2173, 
         nx2175, nx2177, nx2179, nx2181, nx2183, nx2187, nx2189, nx2191, nx2195, 
         nx2203, nx2209, nx2211, nx2213, nx2215, nx2217, nx2219, nx2221, nx2229, 
         nx2231, nx2233, nx2235, nx2237, nx2239, nx2241, nx2245, nx2249, nx2255, 
         nx2257, nx2259, nx2265, nx2269, nx2273, nx2279, nx2281, nx2283, nx2285, 
         nx2291, nx2297, nx2299, nx2301, nx2303, nx2305, nx2307, nx2309, nx2313, 
         nx2317, nx2325, nx2329, nx2335, nx2337, nx2339, nx2341, nx2343, nx2345, 
         nx2347, nx2351, nx2355, nx2359, nx2363, nx2367, nx2373, nx2379, nx2385, 
         nx2387, nx2389, nx2391, nx2393, nx2395, nx2397, nx2401, nx2405, nx2411, 
         nx2413, nx2415, nx2419, nx2423, nx2429, nx2431, nx2433, nx2435, nx2441, 
         nx2445, nx2449, nx2453, nx2459, nx2463, nx2469, nx2475, nx2481, nx2483, 
         nx2485, nx2491, nx2495, nx2499, nx2503, nx2507, nx2511, nx2513, nx2515, 
         nx2519, nx2527, nx2531, nx2535, nx2539, nx2545, nx2549, nx2555, nx2559, 
         nx2565, nx2571, nx2577, nx2579, nx2581, nx2583, nx2585, nx2587, nx2589, 
         nx2597, nx2599, nx2601, nx2603, nx2605, nx2607, nx2609, nx2611, nx2615, 
         nx2617, nx2619, nx2621, nx2625, nx2627, nx2629, nx2631, nx2635, nx2637, 
         nx2639, nx2641, nx2645, nx2647, nx2649, nx2653, nx2661, nx2669, nx2673, 
         nx2679, nx2681, nx2683, nx2689, nx2695, nx2697, nx2699, nx2705, nx2711, 
         nx2713, nx2715, nx2719, nx2723, nx2729, nx2731, nx2733, nx2735, nx2737, 
         nx2739, nx2741, nx2743, nx2747, nx2751, nx2755, nx2759, nx2763, nx2767, 
         nx2771, nx2773, nx2775, nx2779, nx2787, nx2793, nx2795, nx2797, nx2799, 
         nx2801, nx2803, nx2805, nx2813, nx2815, nx2817, nx2819, nx2821, nx2823, 
         nx2825, nx2829, nx2833, nx2841, nx2845, nx2851, nx2853, nx2855, nx2859, 
         nx2863, nx2867, nx2878, nx2886, nx2888, nx2890;
    wire [0:0] \$dummy ;




    nBitRegister_16 RegMultInA (.nBitIn ({A[15],A[14],A[13],A[12],A[11],A[10],
                    A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0]}), .WE (
                    PWR), .Reset (reset), .clk (clk), .Y ({MultA_15,MultA_14,
                    MultA_13,MultA_12,MultA_11,MultA_10,MultA_9,MultA_8,MultA_7,
                    MultA_6,MultA_5,MultA_4,MultA_3,MultA_2,MultA_1,MultA_0})) ;
    nBitRegister_16 RegMultInB (.nBitIn ({B[15],B[14],B[13],B[12],B[11],B[10],
                    B[9],B[8],B[7],B[6],B[5],B[4],B[3],B[2],B[1],B[0]}), .WE (
                    PWR), .Reset (reset), .clk (clk), .Y ({MultB_15,MultB_14,
                    MultB_13,MultB_12,MultB_11,MultB_10,MultB_9,MultB_8,MultB_7,
                    MultB_6,MultB_5,MultB_4,MultB_3,MultB_2,MultB_1,MultB_0})) ;
    nBitRegister_32 RegMultOut (.nBitIn ({Product_31,Product_30,Product_29,
                    Product_28,Product_27,Product_26,Product_25,Product_24,
                    Product_23,Product_22,Product_21,Product_20,Product_19,
                    Product_18,Product_17,Product_16,Product_15,Product_14,
                    Product_13,Product_12,Product_11,Product_10,Product_9,
                    Product_8,Product_7,Product_6,Product_5,Product_4,Product_3,
                    Product_2,Product_1,Product_0}), .WE (PWR), .Reset (reset), 
                    .clk (clk), .Y ({adderB_31,adderB_30,adderB_29,adderB_28,
                    adderB_27,adderB_26,adderB_25,adderB_24,adderB_23,adderB_22,
                    adderB_21,adderB_20,adderB_19,adderB_18,adderB_17,adderB_16,
                    adderB_15,adderB_14,adderB_13,adderB_12,adderB_11,adderB_10,
                    adderB_9,adderB_8,adderB_7,adderB_6,adderB_5,adderB_4,
                    adderB_3,adderB_2,adderB_1,adderB_0})) ;
    nBitRegister_32 BigBoyReg (.nBitIn ({adderOut_31,adderOut_30,adderOut_29,
                    adderOut_28,adderOut_27,adderOut_26,adderOut_25,adderOut_24,
                    adderOut_23,adderOut_22,adderOut_21,adderOut_20,adderOut_19,
                    adderOut_18,adderOut_17,adderOut_16,adderOut_15,adderOut_14,
                    adderOut_13,adderOut_12,adderOut_11,adderOut_10,adderOut_9,
                    adderOut_8,adderOut_7,adderOut_6,adderOut_5,adderOut_4,
                    adderOut_3,adderOut_2,adderOut_1,adderOut_0}), .WE (WE), .Reset (
                    reset), .clk (clk), .Y ({RegOut[31],RegOut[30],RegOut[29],
                    RegOut[28],RegOut[27],RegOut[26],RegOut[25],RegOut[24],
                    RegOut[23],RegOut[22],RegOut[21],RegOut[20],RegOut[19],
                    RegOut[18],RegOut[17],RegOut[16],RegOut[15],RegOut[14],
                    RegOut[13],RegOut[12],RegOut[11],RegOut[10],RegOut[9],
                    RegOut[8],RegOut[7],RegOut[6],RegOut[5],RegOut[4],RegOut[3],
                    RegOut[2],RegOut[1],RegOut[0]})) ;
    full_adder ADD1_generate_adders_0_i_first_adder (.A (RegOut[0]), .B (
               adderB_0), .Cin (MULT1_F_1024), .Sum (adderOut_0), .Cout (
               ADD1_c_array_0)) ;
    full_adder ADD1_generate_adders_1_i_mid_adder (.A (RegOut[1]), .B (adderB_1)
               , .Cin (ADD1_c_array_0), .Sum (adderOut_1), .Cout (ADD1_c_array_1
               )) ;
    full_adder ADD1_generate_adders_2_i_mid_adder (.A (RegOut[2]), .B (adderB_2)
               , .Cin (ADD1_c_array_1), .Sum (adderOut_2), .Cout (ADD1_c_array_2
               )) ;
    full_adder ADD1_generate_adders_3_i_mid_adder (.A (RegOut[3]), .B (adderB_3)
               , .Cin (ADD1_c_array_2), .Sum (adderOut_3), .Cout (ADD1_c_array_3
               )) ;
    full_adder ADD1_generate_adders_4_i_mid_adder (.A (RegOut[4]), .B (adderB_4)
               , .Cin (ADD1_c_array_3), .Sum (adderOut_4), .Cout (ADD1_c_array_4
               )) ;
    full_adder ADD1_generate_adders_5_i_mid_adder (.A (RegOut[5]), .B (adderB_5)
               , .Cin (ADD1_c_array_4), .Sum (adderOut_5), .Cout (ADD1_c_array_5
               )) ;
    full_adder ADD1_generate_adders_6_i_mid_adder (.A (RegOut[6]), .B (adderB_6)
               , .Cin (ADD1_c_array_5), .Sum (adderOut_6), .Cout (ADD1_c_array_6
               )) ;
    full_adder ADD1_generate_adders_7_i_mid_adder (.A (RegOut[7]), .B (adderB_7)
               , .Cin (ADD1_c_array_6), .Sum (adderOut_7), .Cout (ADD1_c_array_7
               )) ;
    full_adder ADD1_generate_adders_8_i_mid_adder (.A (RegOut[8]), .B (adderB_8)
               , .Cin (ADD1_c_array_7), .Sum (adderOut_8), .Cout (ADD1_c_array_8
               )) ;
    full_adder ADD1_generate_adders_9_i_mid_adder (.A (RegOut[9]), .B (adderB_9)
               , .Cin (ADD1_c_array_8), .Sum (adderOut_9), .Cout (ADD1_c_array_9
               )) ;
    full_adder ADD1_generate_adders_10_i_mid_adder (.A (RegOut[10]), .B (
               adderB_10), .Cin (ADD1_c_array_9), .Sum (adderOut_10), .Cout (
               ADD1_c_array_10)) ;
    full_adder ADD1_generate_adders_11_i_mid_adder (.A (RegOut[11]), .B (
               adderB_11), .Cin (ADD1_c_array_10), .Sum (adderOut_11), .Cout (
               ADD1_c_array_11)) ;
    full_adder ADD1_generate_adders_12_i_mid_adder (.A (RegOut[12]), .B (
               adderB_12), .Cin (ADD1_c_array_11), .Sum (adderOut_12), .Cout (
               ADD1_c_array_12)) ;
    full_adder ADD1_generate_adders_13_i_mid_adder (.A (RegOut[13]), .B (
               adderB_13), .Cin (ADD1_c_array_12), .Sum (adderOut_13), .Cout (
               ADD1_c_array_13)) ;
    full_adder ADD1_generate_adders_14_i_mid_adder (.A (RegOut[14]), .B (
               adderB_14), .Cin (ADD1_c_array_13), .Sum (adderOut_14), .Cout (
               ADD1_c_array_14)) ;
    full_adder ADD1_generate_adders_15_i_mid_adder (.A (RegOut[15]), .B (
               adderB_15), .Cin (ADD1_c_array_14), .Sum (adderOut_15), .Cout (
               ADD1_c_array_15)) ;
    full_adder ADD1_generate_adders_16_i_mid_adder (.A (RegOut[16]), .B (
               adderB_16), .Cin (ADD1_c_array_15), .Sum (adderOut_16), .Cout (
               ADD1_c_array_16)) ;
    full_adder ADD1_generate_adders_17_i_mid_adder (.A (RegOut[17]), .B (
               adderB_17), .Cin (ADD1_c_array_16), .Sum (adderOut_17), .Cout (
               ADD1_c_array_17)) ;
    full_adder ADD1_generate_adders_18_i_mid_adder (.A (RegOut[18]), .B (
               adderB_18), .Cin (ADD1_c_array_17), .Sum (adderOut_18), .Cout (
               ADD1_c_array_18)) ;
    full_adder ADD1_generate_adders_19_i_mid_adder (.A (RegOut[19]), .B (
               adderB_19), .Cin (ADD1_c_array_18), .Sum (adderOut_19), .Cout (
               ADD1_c_array_19)) ;
    full_adder ADD1_generate_adders_20_i_mid_adder (.A (RegOut[20]), .B (
               adderB_20), .Cin (ADD1_c_array_19), .Sum (adderOut_20), .Cout (
               ADD1_c_array_20)) ;
    full_adder ADD1_generate_adders_21_i_mid_adder (.A (RegOut[21]), .B (
               adderB_21), .Cin (ADD1_c_array_20), .Sum (adderOut_21), .Cout (
               ADD1_c_array_21)) ;
    full_adder ADD1_generate_adders_22_i_mid_adder (.A (RegOut[22]), .B (
               adderB_22), .Cin (ADD1_c_array_21), .Sum (adderOut_22), .Cout (
               ADD1_c_array_22)) ;
    full_adder ADD1_generate_adders_23_i_mid_adder (.A (RegOut[23]), .B (
               adderB_23), .Cin (ADD1_c_array_22), .Sum (adderOut_23), .Cout (
               ADD1_c_array_23)) ;
    full_adder ADD1_generate_adders_24_i_mid_adder (.A (RegOut[24]), .B (
               adderB_24), .Cin (ADD1_c_array_23), .Sum (adderOut_24), .Cout (
               ADD1_c_array_24)) ;
    full_adder ADD1_generate_adders_25_i_mid_adder (.A (RegOut[25]), .B (
               adderB_25), .Cin (ADD1_c_array_24), .Sum (adderOut_25), .Cout (
               ADD1_c_array_25)) ;
    full_adder ADD1_generate_adders_26_i_mid_adder (.A (RegOut[26]), .B (
               adderB_26), .Cin (ADD1_c_array_25), .Sum (adderOut_26), .Cout (
               ADD1_c_array_26)) ;
    full_adder ADD1_generate_adders_27_i_mid_adder (.A (RegOut[27]), .B (
               adderB_27), .Cin (ADD1_c_array_26), .Sum (adderOut_27), .Cout (
               ADD1_c_array_27)) ;
    full_adder ADD1_generate_adders_28_i_mid_adder (.A (RegOut[28]), .B (
               adderB_28), .Cin (ADD1_c_array_27), .Sum (adderOut_28), .Cout (
               ADD1_c_array_28)) ;
    full_adder ADD1_generate_adders_29_i_mid_adder (.A (RegOut[29]), .B (
               adderB_29), .Cin (ADD1_c_array_28), .Sum (adderOut_29), .Cout (
               ADD1_c_array_29)) ;
    full_adder ADD1_generate_adders_30_i_mid_adder (.A (RegOut[30]), .B (
               adderB_30), .Cin (ADD1_c_array_29), .Sum (adderOut_30), .Cout (
               ADD1_c_array_30)) ;
    full_adder ADD1_generate_adders_31_i_last_adder (.A (RegOut[31]), .B (
               adderB_31), .Cin (ADD1_c_array_30), .Sum (adderOut_31), .Cout (
               \$dummy [0])) ;
    fake_vcc ix458 (.Y (PWR)) ;
    fake_gnd ix456 (.Y (MULT1_F_1024)) ;
    mux21 ix2795 (.Y (Product_15), .A0 (nx497), .A1 (nx2788), .S0 (nx505)) ;
    nand02 ix498 (.Y (nx497), .A0 (MultA_15), .A1 (MultB_0)) ;
    inv01 ix502 (.Y (nx501), .A (MultA_15)) ;
    xnor2 ix506 (.Y (nx505), .A0 (nx1094), .A1 (nx1256)) ;
    nor03 ix1095 (.Y (nx1094), .A0 (nx509), .A1 (nx1495), .A2 (nx2878)) ;
    xnor2 ix510 (.Y (nx509), .A0 (nx938), .A1 (nx1088)) ;
    nor03 ix939 (.Y (nx938), .A0 (nx513), .A1 (nx1363), .A2 (nx2878)) ;
    xnor2 ix514 (.Y (nx513), .A0 (nx794), .A1 (nx932)) ;
    nor03 ix795 (.Y (nx794), .A0 (nx517), .A1 (nx1241), .A2 (nx2878)) ;
    xnor2 ix518 (.Y (nx517), .A0 (nx662), .A1 (nx788)) ;
    nor03 ix663 (.Y (nx662), .A0 (nx521), .A1 (nx1129), .A2 (nx2878)) ;
    xnor2 ix522 (.Y (nx521), .A0 (nx542), .A1 (nx656)) ;
    nor03 ix543 (.Y (nx542), .A0 (nx525), .A1 (nx1027), .A2 (nx2878)) ;
    xnor2 ix526 (.Y (nx525), .A0 (nx434), .A1 (nx536)) ;
    nor03 ix435 (.Y (nx434), .A0 (nx529), .A1 (nx935), .A2 (nx2878)) ;
    xnor2 ix530 (.Y (nx529), .A0 (nx338), .A1 (nx428)) ;
    nor03 ix339 (.Y (nx338), .A0 (nx533), .A1 (nx853), .A2 (nx2878)) ;
    xnor2 ix534 (.Y (nx533), .A0 (nx254), .A1 (nx332)) ;
    nor03 ix255 (.Y (nx254), .A0 (nx537), .A1 (nx781), .A2 (nx2878)) ;
    xnor2 ix538 (.Y (nx537), .A0 (nx182), .A1 (nx248)) ;
    nor03 ix183 (.Y (nx182), .A0 (nx541), .A1 (nx719), .A2 (nx2878)) ;
    xnor2 ix542 (.Y (nx541), .A0 (nx122), .A1 (nx176)) ;
    nor03 ix123 (.Y (nx122), .A0 (nx545), .A1 (nx667), .A2 (nx2878)) ;
    xnor2 ix546 (.Y (nx545), .A0 (nx74), .A1 (nx116)) ;
    nor03 ix75 (.Y (nx74), .A0 (nx549), .A1 (nx625), .A2 (nx2878)) ;
    xnor2 ix550 (.Y (nx549), .A0 (nx38), .A1 (nx68)) ;
    nor03 ix39 (.Y (nx38), .A0 (nx553), .A1 (nx589), .A2 (nx2878)) ;
    xnor2 ix554 (.Y (nx553), .A0 (nx14), .A1 (nx32)) ;
    nor03 ix15 (.Y (nx14), .A0 (nx557), .A1 (nx571), .A2 (nx2878)) ;
    xnor2 ix558 (.Y (nx557), .A0 (nx559), .A1 (nx565)) ;
    nand03 ix560 (.Y (nx559), .A0 (MultA_1), .A1 (MultB_1), .A2 (Product_0)) ;
    xnor2 ix566 (.Y (nx565), .A0 (nx567), .A1 (nx569)) ;
    nand02 ix568 (.Y (nx567), .A0 (MultA_1), .A1 (MultB_1)) ;
    nand02 ix570 (.Y (nx569), .A0 (MultB_2), .A1 (MultA_0)) ;
    inv01 ix572 (.Y (nx571), .A (MultA_2)) ;
    xnor2 ix33 (.Y (nx32), .A0 (nx575), .A1 (nx30)) ;
    nand02 ix576 (.Y (nx575), .A0 (MultA_2), .A1 (MultB_1)) ;
    xnor2 ix31 (.Y (nx30), .A0 (nx22), .A1 (nx583)) ;
    aoi21 ix23 (.Y (nx22), .A0 (nx569), .A1 (nx581), .B0 (nx567)) ;
    nand02 ix582 (.Y (nx581), .A0 (MultB_0), .A1 (MultA_0)) ;
    xnor2 ix584 (.Y (nx583), .A0 (nx585), .A1 (nx587)) ;
    nand02 ix586 (.Y (nx585), .A0 (MultA_1), .A1 (MultB_2)) ;
    nand02 ix588 (.Y (nx587), .A0 (MultB_3), .A1 (MultA_0)) ;
    inv01 ix590 (.Y (nx589), .A (MultA_3)) ;
    xnor2 ix69 (.Y (nx68), .A0 (nx593), .A1 (nx66)) ;
    nand02 ix594 (.Y (nx593), .A0 (MultA_3), .A1 (MultB_1)) ;
    xnor2 ix67 (.Y (nx66), .A0 (nx597), .A1 (nx64)) ;
    aoi32 ix598 (.Y (nx597), .A0 (MultA_2), .A1 (MultB_1), .A2 (nx30), .B0 (nx14
          ), .B1 (nx32)) ;
    xnor2 ix65 (.Y (nx64), .A0 (nx601), .A1 (nx62)) ;
    nand02 ix602 (.Y (nx601), .A0 (MultA_2), .A1 (MultB_2)) ;
    xnor2 ix63 (.Y (nx62), .A0 (nx54), .A1 (nx619)) ;
    oai32 ix55 (.Y (nx54), .A0 (nx607), .A1 (nx609), .A2 (nx587), .B0 (nx611), .B1 (
          nx583)) ;
    inv02 ix608 (.Y (nx607), .A (MultA_1)) ;
    inv01 ix610 (.Y (nx609), .A (MultB_2)) ;
    xnor2 ix620 (.Y (nx619), .A0 (nx621), .A1 (nx623)) ;
    nand02 ix622 (.Y (nx621), .A0 (MultA_1), .A1 (MultB_3)) ;
    nand02 ix624 (.Y (nx623), .A0 (MultB_4), .A1 (MultA_0)) ;
    inv01 ix626 (.Y (nx625), .A (MultA_4)) ;
    xnor2 ix117 (.Y (nx116), .A0 (nx629), .A1 (nx114)) ;
    nand02 ix630 (.Y (nx629), .A0 (MultA_4), .A1 (MultB_1)) ;
    xnor2 ix115 (.Y (nx114), .A0 (nx633), .A1 (nx112)) ;
    aoi32 ix634 (.Y (nx633), .A0 (MultA_3), .A1 (MultB_1), .A2 (nx66), .B0 (nx38
          ), .B1 (nx68)) ;
    xnor2 ix113 (.Y (nx112), .A0 (nx637), .A1 (nx110)) ;
    nand02 ix638 (.Y (nx637), .A0 (MultA_3), .A1 (MultB_2)) ;
    xnor2 ix111 (.Y (nx110), .A0 (nx641), .A1 (nx108)) ;
    aoi32 ix642 (.Y (nx641), .A0 (MultA_2), .A1 (MultB_2), .A2 (nx62), .B0 (nx46
          ), .B1 (nx64)) ;
    xnor2 ix109 (.Y (nx108), .A0 (nx647), .A1 (nx106)) ;
    nand02 ix648 (.Y (nx647), .A0 (MultA_2), .A1 (MultB_3)) ;
    xnor2 ix107 (.Y (nx106), .A0 (nx98), .A1 (nx661)) ;
    oai32 ix99 (.Y (nx98), .A0 (nx607), .A1 (nx653), .A2 (nx623), .B0 (nx655), .B1 (
          nx619)) ;
    inv01 ix654 (.Y (nx653), .A (MultB_3)) ;
    xnor2 ix662 (.Y (nx661), .A0 (nx663), .A1 (nx665)) ;
    nand02 ix664 (.Y (nx663), .A0 (MultA_1), .A1 (MultB_4)) ;
    nand02 ix666 (.Y (nx665), .A0 (MultB_5), .A1 (MultA_0)) ;
    inv01 ix668 (.Y (nx667), .A (MultA_5)) ;
    xnor2 ix177 (.Y (nx176), .A0 (nx671), .A1 (nx174)) ;
    nand02 ix672 (.Y (nx671), .A0 (MultA_5), .A1 (MultB_1)) ;
    xnor2 ix175 (.Y (nx174), .A0 (nx675), .A1 (nx172)) ;
    aoi32 ix676 (.Y (nx675), .A0 (MultA_4), .A1 (MultB_1), .A2 (nx114), .B0 (
          nx74), .B1 (nx116)) ;
    xnor2 ix173 (.Y (nx172), .A0 (nx679), .A1 (nx170)) ;
    nand02 ix680 (.Y (nx679), .A0 (MultA_4), .A1 (MultB_2)) ;
    xnor2 ix171 (.Y (nx170), .A0 (nx683), .A1 (nx168)) ;
    aoi32 ix684 (.Y (nx683), .A0 (MultA_3), .A1 (MultB_2), .A2 (nx110), .B0 (
          nx82), .B1 (nx112)) ;
    xnor2 ix169 (.Y (nx168), .A0 (nx689), .A1 (nx166)) ;
    nand02 ix690 (.Y (nx689), .A0 (MultA_3), .A1 (MultB_3)) ;
    xnor2 ix167 (.Y (nx166), .A0 (nx693), .A1 (nx164)) ;
    aoi32 ix694 (.Y (nx693), .A0 (MultA_2), .A1 (MultB_3), .A2 (nx106), .B0 (
          nx90), .B1 (nx108)) ;
    xnor2 ix165 (.Y (nx164), .A0 (nx699), .A1 (nx162)) ;
    nand02 ix700 (.Y (nx699), .A0 (MultA_2), .A1 (MultB_4)) ;
    xnor2 ix163 (.Y (nx162), .A0 (nx154), .A1 (nx713)) ;
    oai32 ix155 (.Y (nx154), .A0 (nx607), .A1 (nx705), .A2 (nx665), .B0 (nx707)
          , .B1 (nx661)) ;
    inv01 ix706 (.Y (nx705), .A (MultB_4)) ;
    xnor2 ix714 (.Y (nx713), .A0 (nx715), .A1 (nx717)) ;
    nand02 ix716 (.Y (nx715), .A0 (MultA_1), .A1 (MultB_5)) ;
    nand02 ix718 (.Y (nx717), .A0 (MultB_6), .A1 (MultA_0)) ;
    inv01 ix720 (.Y (nx719), .A (MultA_6)) ;
    xnor2 ix249 (.Y (nx248), .A0 (nx723), .A1 (nx246)) ;
    nand02 ix724 (.Y (nx723), .A0 (MultA_6), .A1 (MultB_1)) ;
    xnor2 ix247 (.Y (nx246), .A0 (nx727), .A1 (nx244)) ;
    aoi32 ix728 (.Y (nx727), .A0 (MultA_5), .A1 (MultB_1), .A2 (nx174), .B0 (
          nx122), .B1 (nx176)) ;
    xnor2 ix245 (.Y (nx244), .A0 (nx731), .A1 (nx242)) ;
    nand02 ix732 (.Y (nx731), .A0 (MultA_5), .A1 (MultB_2)) ;
    xnor2 ix243 (.Y (nx242), .A0 (nx735), .A1 (nx240)) ;
    aoi32 ix736 (.Y (nx735), .A0 (MultA_4), .A1 (MultB_2), .A2 (nx170), .B0 (
          nx130), .B1 (nx172)) ;
    xnor2 ix241 (.Y (nx240), .A0 (nx741), .A1 (nx238)) ;
    nand02 ix742 (.Y (nx741), .A0 (MultA_4), .A1 (MultB_3)) ;
    xnor2 ix239 (.Y (nx238), .A0 (nx745), .A1 (nx236)) ;
    aoi32 ix746 (.Y (nx745), .A0 (MultA_3), .A1 (MultB_3), .A2 (nx166), .B0 (
          nx138), .B1 (nx168)) ;
    xnor2 ix237 (.Y (nx236), .A0 (nx751), .A1 (nx234)) ;
    nand02 ix752 (.Y (nx751), .A0 (MultA_3), .A1 (MultB_4)) ;
    xnor2 ix235 (.Y (nx234), .A0 (nx755), .A1 (nx232)) ;
    aoi32 ix756 (.Y (nx755), .A0 (MultA_2), .A1 (MultB_4), .A2 (nx162), .B0 (
          nx146), .B1 (nx164)) ;
    xnor2 ix233 (.Y (nx232), .A0 (nx761), .A1 (nx230)) ;
    nand02 ix762 (.Y (nx761), .A0 (MultA_2), .A1 (MultB_5)) ;
    xnor2 ix231 (.Y (nx230), .A0 (nx222), .A1 (nx775)) ;
    oai32 ix223 (.Y (nx222), .A0 (nx607), .A1 (nx767), .A2 (nx717), .B0 (nx769)
          , .B1 (nx713)) ;
    inv01 ix768 (.Y (nx767), .A (MultB_5)) ;
    xnor2 ix776 (.Y (nx775), .A0 (nx777), .A1 (nx779)) ;
    nand02 ix778 (.Y (nx777), .A0 (MultA_1), .A1 (MultB_6)) ;
    nand02 ix780 (.Y (nx779), .A0 (MultB_7), .A1 (MultA_0)) ;
    inv01 ix782 (.Y (nx781), .A (MultA_7)) ;
    xnor2 ix333 (.Y (nx332), .A0 (nx785), .A1 (nx330)) ;
    nand02 ix786 (.Y (nx785), .A0 (MultA_7), .A1 (MultB_1)) ;
    xnor2 ix331 (.Y (nx330), .A0 (nx789), .A1 (nx328)) ;
    aoi32 ix790 (.Y (nx789), .A0 (MultA_6), .A1 (MultB_1), .A2 (nx246), .B0 (
          nx182), .B1 (nx248)) ;
    xnor2 ix329 (.Y (nx328), .A0 (nx793), .A1 (nx326)) ;
    nand02 ix794 (.Y (nx793), .A0 (MultA_6), .A1 (MultB_2)) ;
    xnor2 ix327 (.Y (nx326), .A0 (nx797), .A1 (nx324)) ;
    aoi32 ix798 (.Y (nx797), .A0 (MultA_5), .A1 (MultB_2), .A2 (nx242), .B0 (
          nx190), .B1 (nx244)) ;
    xnor2 ix325 (.Y (nx324), .A0 (nx803), .A1 (nx322)) ;
    nand02 ix804 (.Y (nx803), .A0 (MultA_5), .A1 (MultB_3)) ;
    xnor2 ix323 (.Y (nx322), .A0 (nx807), .A1 (nx320)) ;
    aoi32 ix808 (.Y (nx807), .A0 (MultA_4), .A1 (MultB_3), .A2 (nx238), .B0 (
          nx198), .B1 (nx240)) ;
    xnor2 ix321 (.Y (nx320), .A0 (nx813), .A1 (nx318)) ;
    nand02 ix814 (.Y (nx813), .A0 (MultA_4), .A1 (MultB_4)) ;
    xnor2 ix319 (.Y (nx318), .A0 (nx817), .A1 (nx316)) ;
    aoi32 ix818 (.Y (nx817), .A0 (MultA_3), .A1 (MultB_4), .A2 (nx234), .B0 (
          nx206), .B1 (nx236)) ;
    xnor2 ix317 (.Y (nx316), .A0 (nx823), .A1 (nx314)) ;
    nand02 ix824 (.Y (nx823), .A0 (MultA_3), .A1 (MultB_5)) ;
    xnor2 ix315 (.Y (nx314), .A0 (nx827), .A1 (nx312)) ;
    aoi32 ix828 (.Y (nx827), .A0 (MultA_2), .A1 (MultB_5), .A2 (nx230), .B0 (
          nx214), .B1 (nx232)) ;
    xnor2 ix313 (.Y (nx312), .A0 (nx833), .A1 (nx310)) ;
    nand02 ix834 (.Y (nx833), .A0 (MultA_2), .A1 (MultB_6)) ;
    xnor2 ix311 (.Y (nx310), .A0 (nx302), .A1 (nx847)) ;
    oai32 ix303 (.Y (nx302), .A0 (nx607), .A1 (nx839), .A2 (nx779), .B0 (nx841)
          , .B1 (nx775)) ;
    inv01 ix840 (.Y (nx839), .A (MultB_6)) ;
    xnor2 ix848 (.Y (nx847), .A0 (nx849), .A1 (nx851)) ;
    nand02 ix850 (.Y (nx849), .A0 (MultA_1), .A1 (MultB_7)) ;
    nand02 ix852 (.Y (nx851), .A0 (MultB_8), .A1 (MultA_0)) ;
    inv01 ix854 (.Y (nx853), .A (MultA_8)) ;
    xnor2 ix429 (.Y (nx428), .A0 (nx857), .A1 (nx426)) ;
    nand02 ix858 (.Y (nx857), .A0 (MultA_8), .A1 (MultB_1)) ;
    xnor2 ix427 (.Y (nx426), .A0 (nx861), .A1 (nx424)) ;
    aoi32 ix862 (.Y (nx861), .A0 (MultA_7), .A1 (MultB_1), .A2 (nx330), .B0 (
          nx254), .B1 (nx332)) ;
    xnor2 ix425 (.Y (nx424), .A0 (nx865), .A1 (nx422)) ;
    nand02 ix866 (.Y (nx865), .A0 (MultA_7), .A1 (MultB_2)) ;
    xnor2 ix423 (.Y (nx422), .A0 (nx869), .A1 (nx420)) ;
    aoi32 ix870 (.Y (nx869), .A0 (MultA_6), .A1 (MultB_2), .A2 (nx326), .B0 (
          nx262), .B1 (nx328)) ;
    xnor2 ix421 (.Y (nx420), .A0 (nx875), .A1 (nx418)) ;
    nand02 ix876 (.Y (nx875), .A0 (MultA_6), .A1 (MultB_3)) ;
    xnor2 ix419 (.Y (nx418), .A0 (nx879), .A1 (nx416)) ;
    aoi32 ix880 (.Y (nx879), .A0 (MultA_5), .A1 (MultB_3), .A2 (nx322), .B0 (
          nx270), .B1 (nx324)) ;
    xnor2 ix417 (.Y (nx416), .A0 (nx885), .A1 (nx414)) ;
    nand02 ix886 (.Y (nx885), .A0 (MultA_5), .A1 (MultB_4)) ;
    xnor2 ix415 (.Y (nx414), .A0 (nx889), .A1 (nx412)) ;
    aoi32 ix890 (.Y (nx889), .A0 (MultA_4), .A1 (MultB_4), .A2 (nx318), .B0 (
          nx278), .B1 (nx320)) ;
    xnor2 ix413 (.Y (nx412), .A0 (nx895), .A1 (nx410)) ;
    nand02 ix896 (.Y (nx895), .A0 (MultA_4), .A1 (MultB_5)) ;
    xnor2 ix411 (.Y (nx410), .A0 (nx899), .A1 (nx408)) ;
    aoi32 ix900 (.Y (nx899), .A0 (MultA_3), .A1 (MultB_5), .A2 (nx314), .B0 (
          nx286), .B1 (nx316)) ;
    xnor2 ix409 (.Y (nx408), .A0 (nx905), .A1 (nx406)) ;
    nand02 ix906 (.Y (nx905), .A0 (MultA_3), .A1 (MultB_6)) ;
    xnor2 ix407 (.Y (nx406), .A0 (nx909), .A1 (nx404)) ;
    aoi32 ix910 (.Y (nx909), .A0 (MultA_2), .A1 (MultB_6), .A2 (nx310), .B0 (
          nx294), .B1 (nx312)) ;
    xnor2 ix405 (.Y (nx404), .A0 (nx915), .A1 (nx402)) ;
    nand02 ix916 (.Y (nx915), .A0 (MultA_2), .A1 (MultB_7)) ;
    xnor2 ix403 (.Y (nx402), .A0 (nx394), .A1 (nx929)) ;
    oai32 ix395 (.Y (nx394), .A0 (nx607), .A1 (nx921), .A2 (nx851), .B0 (nx923)
          , .B1 (nx847)) ;
    inv01 ix922 (.Y (nx921), .A (MultB_7)) ;
    xnor2 ix930 (.Y (nx929), .A0 (nx931), .A1 (nx933)) ;
    nand02 ix932 (.Y (nx931), .A0 (MultA_1), .A1 (MultB_8)) ;
    nand02 ix934 (.Y (nx933), .A0 (MultB_9), .A1 (MultA_0)) ;
    inv01 ix936 (.Y (nx935), .A (MultA_9)) ;
    xnor2 ix537 (.Y (nx536), .A0 (nx939), .A1 (nx534)) ;
    nand02 ix940 (.Y (nx939), .A0 (MultA_9), .A1 (MultB_1)) ;
    xnor2 ix535 (.Y (nx534), .A0 (nx943), .A1 (nx532)) ;
    aoi32 ix944 (.Y (nx943), .A0 (MultA_8), .A1 (MultB_1), .A2 (nx426), .B0 (
          nx338), .B1 (nx428)) ;
    xnor2 ix533 (.Y (nx532), .A0 (nx947), .A1 (nx530)) ;
    nand02 ix948 (.Y (nx947), .A0 (MultA_8), .A1 (MultB_2)) ;
    xnor2 ix531 (.Y (nx530), .A0 (nx951), .A1 (nx528)) ;
    aoi32 ix952 (.Y (nx951), .A0 (MultA_7), .A1 (MultB_2), .A2 (nx422), .B0 (
          nx346), .B1 (nx424)) ;
    xnor2 ix529 (.Y (nx528), .A0 (nx957), .A1 (nx526)) ;
    nand02 ix958 (.Y (nx957), .A0 (MultA_7), .A1 (MultB_3)) ;
    xnor2 ix527 (.Y (nx526), .A0 (nx961), .A1 (nx524)) ;
    aoi32 ix962 (.Y (nx961), .A0 (MultA_6), .A1 (MultB_3), .A2 (nx418), .B0 (
          nx354), .B1 (nx420)) ;
    xnor2 ix525 (.Y (nx524), .A0 (nx967), .A1 (nx522)) ;
    nand02 ix968 (.Y (nx967), .A0 (MultA_6), .A1 (MultB_4)) ;
    xnor2 ix523 (.Y (nx522), .A0 (nx971), .A1 (nx520)) ;
    aoi32 ix972 (.Y (nx971), .A0 (MultA_5), .A1 (MultB_4), .A2 (nx414), .B0 (
          nx362), .B1 (nx416)) ;
    xnor2 ix521 (.Y (nx520), .A0 (nx977), .A1 (nx518)) ;
    nand02 ix978 (.Y (nx977), .A0 (MultA_5), .A1 (MultB_5)) ;
    xnor2 ix519 (.Y (nx518), .A0 (nx981), .A1 (nx516)) ;
    aoi32 ix982 (.Y (nx981), .A0 (MultA_4), .A1 (MultB_5), .A2 (nx410), .B0 (
          nx370), .B1 (nx412)) ;
    xnor2 ix517 (.Y (nx516), .A0 (nx987), .A1 (nx514)) ;
    nand02 ix988 (.Y (nx987), .A0 (MultA_4), .A1 (MultB_6)) ;
    xnor2 ix515 (.Y (nx514), .A0 (nx991), .A1 (nx512)) ;
    aoi32 ix992 (.Y (nx991), .A0 (MultA_3), .A1 (MultB_6), .A2 (nx406), .B0 (
          nx378), .B1 (nx408)) ;
    xnor2 ix513 (.Y (nx512), .A0 (nx997), .A1 (nx510)) ;
    nand02 ix998 (.Y (nx997), .A0 (MultA_3), .A1 (MultB_7)) ;
    xnor2 ix511 (.Y (nx510), .A0 (nx1001), .A1 (nx508)) ;
    aoi32 ix1002 (.Y (nx1001), .A0 (MultA_2), .A1 (MultB_7), .A2 (nx402), .B0 (
          nx386), .B1 (nx404)) ;
    xnor2 ix509 (.Y (nx508), .A0 (nx1007), .A1 (nx506)) ;
    nand02 ix1008 (.Y (nx1007), .A0 (MultA_2), .A1 (MultB_8)) ;
    xnor2 ix507 (.Y (nx506), .A0 (nx498), .A1 (nx1021)) ;
    oai32 ix499 (.Y (nx498), .A0 (nx607), .A1 (nx1013), .A2 (nx933), .B0 (nx1015
          ), .B1 (nx929)) ;
    inv01 ix1014 (.Y (nx1013), .A (MultB_8)) ;
    xnor2 ix1022 (.Y (nx1021), .A0 (nx1023), .A1 (nx1025)) ;
    nand02 ix1024 (.Y (nx1023), .A0 (MultA_1), .A1 (MultB_9)) ;
    nand02 ix1026 (.Y (nx1025), .A0 (MultB_10), .A1 (MultA_0)) ;
    inv01 ix1028 (.Y (nx1027), .A (MultA_10)) ;
    xnor2 ix657 (.Y (nx656), .A0 (nx1031), .A1 (nx654)) ;
    nand02 ix1032 (.Y (nx1031), .A0 (MultA_10), .A1 (MultB_1)) ;
    xnor2 ix655 (.Y (nx654), .A0 (nx1035), .A1 (nx652)) ;
    aoi32 ix1036 (.Y (nx1035), .A0 (MultA_9), .A1 (MultB_1), .A2 (nx534), .B0 (
          nx434), .B1 (nx536)) ;
    xnor2 ix653 (.Y (nx652), .A0 (nx1039), .A1 (nx650)) ;
    nand02 ix1040 (.Y (nx1039), .A0 (MultA_9), .A1 (MultB_2)) ;
    xnor2 ix651 (.Y (nx650), .A0 (nx1043), .A1 (nx648)) ;
    aoi32 ix1044 (.Y (nx1043), .A0 (MultA_8), .A1 (MultB_2), .A2 (nx530), .B0 (
          nx442), .B1 (nx532)) ;
    xnor2 ix649 (.Y (nx648), .A0 (nx1049), .A1 (nx646)) ;
    nand02 ix1050 (.Y (nx1049), .A0 (MultA_8), .A1 (MultB_3)) ;
    xnor2 ix647 (.Y (nx646), .A0 (nx1053), .A1 (nx644)) ;
    aoi32 ix1054 (.Y (nx1053), .A0 (MultA_7), .A1 (MultB_3), .A2 (nx526), .B0 (
          nx450), .B1 (nx528)) ;
    xnor2 ix645 (.Y (nx644), .A0 (nx1059), .A1 (nx642)) ;
    nand02 ix1060 (.Y (nx1059), .A0 (MultA_7), .A1 (MultB_4)) ;
    xnor2 ix643 (.Y (nx642), .A0 (nx1063), .A1 (nx640)) ;
    aoi32 ix1064 (.Y (nx1063), .A0 (MultA_6), .A1 (MultB_4), .A2 (nx522), .B0 (
          nx458), .B1 (nx524)) ;
    xnor2 ix641 (.Y (nx640), .A0 (nx1069), .A1 (nx638)) ;
    nand02 ix1070 (.Y (nx1069), .A0 (MultA_6), .A1 (MultB_5)) ;
    xnor2 ix639 (.Y (nx638), .A0 (nx1073), .A1 (nx636)) ;
    aoi32 ix1074 (.Y (nx1073), .A0 (MultA_5), .A1 (MultB_5), .A2 (nx518), .B0 (
          nx466), .B1 (nx520)) ;
    xnor2 ix637 (.Y (nx636), .A0 (nx1079), .A1 (nx634)) ;
    nand02 ix1080 (.Y (nx1079), .A0 (MultA_5), .A1 (MultB_6)) ;
    xnor2 ix635 (.Y (nx634), .A0 (nx1083), .A1 (nx632)) ;
    aoi32 ix1084 (.Y (nx1083), .A0 (MultA_4), .A1 (MultB_6), .A2 (nx514), .B0 (
          nx474), .B1 (nx516)) ;
    xnor2 ix633 (.Y (nx632), .A0 (nx1089), .A1 (nx630)) ;
    nand02 ix1090 (.Y (nx1089), .A0 (MultA_4), .A1 (MultB_7)) ;
    xnor2 ix631 (.Y (nx630), .A0 (nx1093), .A1 (nx628)) ;
    aoi32 ix1094 (.Y (nx1093), .A0 (MultA_3), .A1 (MultB_7), .A2 (nx510), .B0 (
          nx482), .B1 (nx512)) ;
    xnor2 ix629 (.Y (nx628), .A0 (nx1099), .A1 (nx626)) ;
    nand02 ix1100 (.Y (nx1099), .A0 (MultA_3), .A1 (MultB_8)) ;
    xnor2 ix627 (.Y (nx626), .A0 (nx1103), .A1 (nx624)) ;
    aoi32 ix1104 (.Y (nx1103), .A0 (MultA_2), .A1 (MultB_8), .A2 (nx506), .B0 (
          nx490), .B1 (nx508)) ;
    xnor2 ix625 (.Y (nx624), .A0 (nx1109), .A1 (nx622)) ;
    nand02 ix1110 (.Y (nx1109), .A0 (MultA_2), .A1 (MultB_9)) ;
    xnor2 ix623 (.Y (nx622), .A0 (nx614), .A1 (nx1123)) ;
    oai32 ix615 (.Y (nx614), .A0 (nx607), .A1 (nx1115), .A2 (nx1025), .B0 (
          nx1117), .B1 (nx1021)) ;
    inv01 ix1116 (.Y (nx1115), .A (MultB_9)) ;
    xnor2 ix1124 (.Y (nx1123), .A0 (nx1125), .A1 (nx1127)) ;
    nand02 ix1126 (.Y (nx1125), .A0 (MultA_1), .A1 (MultB_10)) ;
    nand02 ix1128 (.Y (nx1127), .A0 (MultB_11), .A1 (MultA_0)) ;
    inv01 ix1130 (.Y (nx1129), .A (MultA_11)) ;
    xnor2 ix789 (.Y (nx788), .A0 (nx1133), .A1 (nx786)) ;
    nand02 ix1134 (.Y (nx1133), .A0 (MultA_11), .A1 (MultB_1)) ;
    xnor2 ix787 (.Y (nx786), .A0 (nx1137), .A1 (nx784)) ;
    aoi32 ix1138 (.Y (nx1137), .A0 (MultA_10), .A1 (MultB_1), .A2 (nx654), .B0 (
          nx542), .B1 (nx656)) ;
    xnor2 ix785 (.Y (nx784), .A0 (nx1141), .A1 (nx782)) ;
    nand02 ix1142 (.Y (nx1141), .A0 (MultA_10), .A1 (MultB_2)) ;
    xnor2 ix783 (.Y (nx782), .A0 (nx1145), .A1 (nx780)) ;
    aoi32 ix1146 (.Y (nx1145), .A0 (MultA_9), .A1 (MultB_2), .A2 (nx650), .B0 (
          nx550), .B1 (nx652)) ;
    xnor2 ix781 (.Y (nx780), .A0 (nx1151), .A1 (nx778)) ;
    nand02 ix1152 (.Y (nx1151), .A0 (MultA_9), .A1 (MultB_3)) ;
    xnor2 ix779 (.Y (nx778), .A0 (nx1155), .A1 (nx776)) ;
    aoi32 ix1156 (.Y (nx1155), .A0 (MultA_8), .A1 (MultB_3), .A2 (nx646), .B0 (
          nx558), .B1 (nx648)) ;
    xnor2 ix777 (.Y (nx776), .A0 (nx1161), .A1 (nx774)) ;
    nand02 ix1162 (.Y (nx1161), .A0 (MultA_8), .A1 (MultB_4)) ;
    xnor2 ix775 (.Y (nx774), .A0 (nx1165), .A1 (nx772)) ;
    aoi32 ix1166 (.Y (nx1165), .A0 (MultA_7), .A1 (MultB_4), .A2 (nx642), .B0 (
          nx566), .B1 (nx644)) ;
    xnor2 ix773 (.Y (nx772), .A0 (nx1171), .A1 (nx770)) ;
    nand02 ix1172 (.Y (nx1171), .A0 (MultA_7), .A1 (MultB_5)) ;
    xnor2 ix771 (.Y (nx770), .A0 (nx1175), .A1 (nx768)) ;
    aoi32 ix1176 (.Y (nx1175), .A0 (MultA_6), .A1 (MultB_5), .A2 (nx638), .B0 (
          nx574), .B1 (nx640)) ;
    xnor2 ix769 (.Y (nx768), .A0 (nx1181), .A1 (nx766)) ;
    nand02 ix1182 (.Y (nx1181), .A0 (MultA_6), .A1 (MultB_6)) ;
    xnor2 ix767 (.Y (nx766), .A0 (nx1185), .A1 (nx764)) ;
    aoi32 ix1186 (.Y (nx1185), .A0 (MultA_5), .A1 (MultB_6), .A2 (nx634), .B0 (
          nx582), .B1 (nx636)) ;
    xnor2 ix765 (.Y (nx764), .A0 (nx1191), .A1 (nx762)) ;
    nand02 ix1192 (.Y (nx1191), .A0 (MultA_5), .A1 (MultB_7)) ;
    xnor2 ix763 (.Y (nx762), .A0 (nx1195), .A1 (nx760)) ;
    aoi32 ix1196 (.Y (nx1195), .A0 (MultA_4), .A1 (MultB_7), .A2 (nx630), .B0 (
          nx590), .B1 (nx632)) ;
    xnor2 ix761 (.Y (nx760), .A0 (nx1201), .A1 (nx758)) ;
    nand02 ix1202 (.Y (nx1201), .A0 (MultA_4), .A1 (MultB_8)) ;
    xnor2 ix759 (.Y (nx758), .A0 (nx1205), .A1 (nx756)) ;
    aoi32 ix1206 (.Y (nx1205), .A0 (MultA_3), .A1 (MultB_8), .A2 (nx626), .B0 (
          nx598), .B1 (nx628)) ;
    xnor2 ix757 (.Y (nx756), .A0 (nx1211), .A1 (nx754)) ;
    nand02 ix1212 (.Y (nx1211), .A0 (MultA_3), .A1 (MultB_9)) ;
    xnor2 ix755 (.Y (nx754), .A0 (nx1215), .A1 (nx752)) ;
    aoi32 ix1216 (.Y (nx1215), .A0 (MultA_2), .A1 (MultB_9), .A2 (nx622), .B0 (
          nx606), .B1 (nx624)) ;
    xnor2 ix753 (.Y (nx752), .A0 (nx1221), .A1 (nx750)) ;
    nand02 ix1222 (.Y (nx1221), .A0 (MultA_2), .A1 (MultB_10)) ;
    xnor2 ix751 (.Y (nx750), .A0 (nx742), .A1 (nx1235)) ;
    oai32 ix743 (.Y (nx742), .A0 (nx607), .A1 (nx1227), .A2 (nx1127), .B0 (
          nx1229), .B1 (nx1123)) ;
    inv01 ix1228 (.Y (nx1227), .A (MultB_10)) ;
    xnor2 ix1236 (.Y (nx1235), .A0 (nx1237), .A1 (nx1239)) ;
    nand02 ix1238 (.Y (nx1237), .A0 (MultA_1), .A1 (MultB_11)) ;
    nand02 ix1240 (.Y (nx1239), .A0 (MultB_12), .A1 (MultA_0)) ;
    inv01 ix1242 (.Y (nx1241), .A (MultA_12)) ;
    xnor2 ix933 (.Y (nx932), .A0 (nx1245), .A1 (nx930)) ;
    nand02 ix1246 (.Y (nx1245), .A0 (MultA_12), .A1 (MultB_1)) ;
    xnor2 ix931 (.Y (nx930), .A0 (nx1249), .A1 (nx928)) ;
    aoi32 ix1250 (.Y (nx1249), .A0 (MultA_11), .A1 (MultB_1), .A2 (nx786), .B0 (
          nx662), .B1 (nx788)) ;
    xnor2 ix929 (.Y (nx928), .A0 (nx1253), .A1 (nx926)) ;
    nand02 ix1254 (.Y (nx1253), .A0 (MultA_11), .A1 (MultB_2)) ;
    xnor2 ix927 (.Y (nx926), .A0 (nx1257), .A1 (nx924)) ;
    aoi32 ix1258 (.Y (nx1257), .A0 (MultA_10), .A1 (MultB_2), .A2 (nx782), .B0 (
          nx670), .B1 (nx784)) ;
    xnor2 ix925 (.Y (nx924), .A0 (nx1263), .A1 (nx922)) ;
    nand02 ix1264 (.Y (nx1263), .A0 (MultA_10), .A1 (MultB_3)) ;
    xnor2 ix923 (.Y (nx922), .A0 (nx1267), .A1 (nx920)) ;
    aoi32 ix1268 (.Y (nx1267), .A0 (MultA_9), .A1 (MultB_3), .A2 (nx778), .B0 (
          nx678), .B1 (nx780)) ;
    xnor2 ix921 (.Y (nx920), .A0 (nx1273), .A1 (nx918)) ;
    nand02 ix1274 (.Y (nx1273), .A0 (MultA_9), .A1 (MultB_4)) ;
    xnor2 ix919 (.Y (nx918), .A0 (nx1277), .A1 (nx916)) ;
    aoi32 ix1278 (.Y (nx1277), .A0 (MultA_8), .A1 (MultB_4), .A2 (nx774), .B0 (
          nx686), .B1 (nx776)) ;
    xnor2 ix917 (.Y (nx916), .A0 (nx1283), .A1 (nx914)) ;
    nand02 ix1284 (.Y (nx1283), .A0 (MultA_8), .A1 (MultB_5)) ;
    xnor2 ix915 (.Y (nx914), .A0 (nx1287), .A1 (nx912)) ;
    aoi32 ix1288 (.Y (nx1287), .A0 (MultA_7), .A1 (MultB_5), .A2 (nx770), .B0 (
          nx694), .B1 (nx772)) ;
    xnor2 ix913 (.Y (nx912), .A0 (nx1293), .A1 (nx910)) ;
    nand02 ix1294 (.Y (nx1293), .A0 (MultA_7), .A1 (MultB_6)) ;
    xnor2 ix911 (.Y (nx910), .A0 (nx1297), .A1 (nx908)) ;
    aoi32 ix1298 (.Y (nx1297), .A0 (MultA_6), .A1 (MultB_6), .A2 (nx766), .B0 (
          nx702), .B1 (nx768)) ;
    xnor2 ix909 (.Y (nx908), .A0 (nx1303), .A1 (nx906)) ;
    nand02 ix1304 (.Y (nx1303), .A0 (MultA_6), .A1 (MultB_7)) ;
    xnor2 ix907 (.Y (nx906), .A0 (nx1307), .A1 (nx904)) ;
    aoi32 ix1308 (.Y (nx1307), .A0 (MultA_5), .A1 (MultB_7), .A2 (nx762), .B0 (
          nx710), .B1 (nx764)) ;
    xnor2 ix905 (.Y (nx904), .A0 (nx1313), .A1 (nx902)) ;
    nand02 ix1314 (.Y (nx1313), .A0 (MultA_5), .A1 (MultB_8)) ;
    xnor2 ix903 (.Y (nx902), .A0 (nx1317), .A1 (nx900)) ;
    aoi32 ix1318 (.Y (nx1317), .A0 (MultA_4), .A1 (MultB_8), .A2 (nx758), .B0 (
          nx718), .B1 (nx760)) ;
    xnor2 ix901 (.Y (nx900), .A0 (nx1323), .A1 (nx898)) ;
    nand02 ix1324 (.Y (nx1323), .A0 (MultA_4), .A1 (MultB_9)) ;
    xnor2 ix899 (.Y (nx898), .A0 (nx1327), .A1 (nx896)) ;
    aoi32 ix1328 (.Y (nx1327), .A0 (MultA_3), .A1 (MultB_9), .A2 (nx754), .B0 (
          nx726), .B1 (nx756)) ;
    xnor2 ix897 (.Y (nx896), .A0 (nx1333), .A1 (nx894)) ;
    nand02 ix1334 (.Y (nx1333), .A0 (MultA_3), .A1 (MultB_10)) ;
    xnor2 ix895 (.Y (nx894), .A0 (nx1337), .A1 (nx892)) ;
    aoi32 ix1338 (.Y (nx1337), .A0 (MultA_2), .A1 (MultB_10), .A2 (nx750), .B0 (
          nx734), .B1 (nx752)) ;
    xnor2 ix893 (.Y (nx892), .A0 (nx1343), .A1 (nx890)) ;
    nand02 ix1344 (.Y (nx1343), .A0 (MultA_2), .A1 (MultB_11)) ;
    xnor2 ix891 (.Y (nx890), .A0 (nx882), .A1 (nx1357)) ;
    oai32 ix883 (.Y (nx882), .A0 (nx607), .A1 (nx1349), .A2 (nx1239), .B0 (
          nx1351), .B1 (nx1235)) ;
    inv01 ix1350 (.Y (nx1349), .A (MultB_11)) ;
    xnor2 ix1358 (.Y (nx1357), .A0 (nx1359), .A1 (nx1361)) ;
    nand02 ix1360 (.Y (nx1359), .A0 (MultA_1), .A1 (MultB_12)) ;
    nand02 ix1362 (.Y (nx1361), .A0 (MultB_13), .A1 (MultA_0)) ;
    inv01 ix1364 (.Y (nx1363), .A (MultA_13)) ;
    xnor2 ix1089 (.Y (nx1088), .A0 (nx1367), .A1 (nx1086)) ;
    nand02 ix1368 (.Y (nx1367), .A0 (MultA_13), .A1 (MultB_1)) ;
    xnor2 ix1087 (.Y (nx1086), .A0 (nx1371), .A1 (nx1084)) ;
    aoi32 ix1372 (.Y (nx1371), .A0 (MultA_12), .A1 (MultB_1), .A2 (nx930), .B0 (
          nx794), .B1 (nx932)) ;
    xnor2 ix1085 (.Y (nx1084), .A0 (nx1375), .A1 (nx1082)) ;
    nand02 ix1376 (.Y (nx1375), .A0 (MultA_12), .A1 (MultB_2)) ;
    xnor2 ix1083 (.Y (nx1082), .A0 (nx1379), .A1 (nx1080)) ;
    aoi32 ix1380 (.Y (nx1379), .A0 (MultA_11), .A1 (MultB_2), .A2 (nx926), .B0 (
          nx802), .B1 (nx928)) ;
    xnor2 ix1081 (.Y (nx1080), .A0 (nx1385), .A1 (nx1078)) ;
    nand02 ix1386 (.Y (nx1385), .A0 (MultA_11), .A1 (MultB_3)) ;
    xnor2 ix1079 (.Y (nx1078), .A0 (nx1389), .A1 (nx1076)) ;
    aoi32 ix1390 (.Y (nx1389), .A0 (MultA_10), .A1 (MultB_3), .A2 (nx922), .B0 (
          nx810), .B1 (nx924)) ;
    xnor2 ix1077 (.Y (nx1076), .A0 (nx1395), .A1 (nx1074)) ;
    nand02 ix1396 (.Y (nx1395), .A0 (MultA_10), .A1 (MultB_4)) ;
    xnor2 ix1075 (.Y (nx1074), .A0 (nx1399), .A1 (nx1072)) ;
    aoi32 ix1400 (.Y (nx1399), .A0 (MultA_9), .A1 (MultB_4), .A2 (nx918), .B0 (
          nx818), .B1 (nx920)) ;
    xnor2 ix1073 (.Y (nx1072), .A0 (nx1405), .A1 (nx1070)) ;
    nand02 ix1406 (.Y (nx1405), .A0 (MultA_9), .A1 (MultB_5)) ;
    xnor2 ix1071 (.Y (nx1070), .A0 (nx1409), .A1 (nx1068)) ;
    aoi32 ix1410 (.Y (nx1409), .A0 (MultA_8), .A1 (MultB_5), .A2 (nx914), .B0 (
          nx826), .B1 (nx916)) ;
    xnor2 ix1069 (.Y (nx1068), .A0 (nx1415), .A1 (nx1066)) ;
    nand02 ix1416 (.Y (nx1415), .A0 (MultA_8), .A1 (MultB_6)) ;
    xnor2 ix1067 (.Y (nx1066), .A0 (nx1419), .A1 (nx1064)) ;
    aoi32 ix1420 (.Y (nx1419), .A0 (MultA_7), .A1 (MultB_6), .A2 (nx910), .B0 (
          nx834), .B1 (nx912)) ;
    xnor2 ix1065 (.Y (nx1064), .A0 (nx1425), .A1 (nx1062)) ;
    nand02 ix1426 (.Y (nx1425), .A0 (MultA_7), .A1 (MultB_7)) ;
    xnor2 ix1063 (.Y (nx1062), .A0 (nx1429), .A1 (nx1060)) ;
    aoi32 ix1430 (.Y (nx1429), .A0 (MultA_6), .A1 (MultB_7), .A2 (nx906), .B0 (
          nx842), .B1 (nx908)) ;
    xnor2 ix1061 (.Y (nx1060), .A0 (nx1435), .A1 (nx1058)) ;
    nand02 ix1436 (.Y (nx1435), .A0 (MultA_6), .A1 (MultB_8)) ;
    xnor2 ix1059 (.Y (nx1058), .A0 (nx1439), .A1 (nx1056)) ;
    aoi32 ix1440 (.Y (nx1439), .A0 (MultA_5), .A1 (MultB_8), .A2 (nx902), .B0 (
          nx850), .B1 (nx904)) ;
    xnor2 ix1057 (.Y (nx1056), .A0 (nx1445), .A1 (nx1054)) ;
    nand02 ix1446 (.Y (nx1445), .A0 (MultA_5), .A1 (MultB_9)) ;
    xnor2 ix1055 (.Y (nx1054), .A0 (nx1449), .A1 (nx1052)) ;
    aoi32 ix1450 (.Y (nx1449), .A0 (MultA_4), .A1 (MultB_9), .A2 (nx898), .B0 (
          nx858), .B1 (nx900)) ;
    xnor2 ix1053 (.Y (nx1052), .A0 (nx1455), .A1 (nx1050)) ;
    nand02 ix1456 (.Y (nx1455), .A0 (MultA_4), .A1 (MultB_10)) ;
    xnor2 ix1051 (.Y (nx1050), .A0 (nx1459), .A1 (nx1048)) ;
    aoi32 ix1460 (.Y (nx1459), .A0 (MultA_3), .A1 (MultB_10), .A2 (nx894), .B0 (
          nx866), .B1 (nx896)) ;
    xnor2 ix1049 (.Y (nx1048), .A0 (nx1465), .A1 (nx1046)) ;
    nand02 ix1466 (.Y (nx1465), .A0 (MultA_3), .A1 (MultB_11)) ;
    xnor2 ix1047 (.Y (nx1046), .A0 (nx1469), .A1 (nx1044)) ;
    aoi32 ix1470 (.Y (nx1469), .A0 (MultA_2), .A1 (MultB_11), .A2 (nx890), .B0 (
          nx874), .B1 (nx892)) ;
    xnor2 ix1045 (.Y (nx1044), .A0 (nx1475), .A1 (nx1042)) ;
    nand02 ix1476 (.Y (nx1475), .A0 (MultA_2), .A1 (MultB_12)) ;
    xnor2 ix1043 (.Y (nx1042), .A0 (nx1034), .A1 (nx1489)) ;
    oai32 ix1035 (.Y (nx1034), .A0 (nx607), .A1 (nx1481), .A2 (nx1361), .B0 (
          nx1483), .B1 (nx1357)) ;
    inv01 ix1482 (.Y (nx1481), .A (MultB_12)) ;
    xnor2 ix1490 (.Y (nx1489), .A0 (nx1491), .A1 (nx1493)) ;
    nand02 ix1492 (.Y (nx1491), .A0 (MultA_1), .A1 (MultB_13)) ;
    nand02 ix1494 (.Y (nx1493), .A0 (MultB_14), .A1 (MultA_0)) ;
    inv01 ix1496 (.Y (nx1495), .A (MultA_14)) ;
    xnor2 ix1257 (.Y (nx1256), .A0 (nx1499), .A1 (nx1254)) ;
    nand02 ix1500 (.Y (nx1499), .A0 (MultA_14), .A1 (MultB_1)) ;
    xnor2 ix1255 (.Y (nx1254), .A0 (nx1503), .A1 (nx1252)) ;
    aoi32 ix1504 (.Y (nx1503), .A0 (MultA_13), .A1 (MultB_1), .A2 (nx1086), .B0 (
          nx938), .B1 (nx1088)) ;
    xnor2 ix1253 (.Y (nx1252), .A0 (nx1507), .A1 (nx1250)) ;
    nand02 ix1508 (.Y (nx1507), .A0 (MultA_13), .A1 (MultB_2)) ;
    xnor2 ix1251 (.Y (nx1250), .A0 (nx1511), .A1 (nx1248)) ;
    aoi32 ix1512 (.Y (nx1511), .A0 (MultA_12), .A1 (MultB_2), .A2 (nx1082), .B0 (
          nx946), .B1 (nx1084)) ;
    xnor2 ix1249 (.Y (nx1248), .A0 (nx1517), .A1 (nx1246)) ;
    nand02 ix1518 (.Y (nx1517), .A0 (MultA_12), .A1 (MultB_3)) ;
    xnor2 ix1247 (.Y (nx1246), .A0 (nx1521), .A1 (nx1244)) ;
    aoi32 ix1522 (.Y (nx1521), .A0 (MultA_11), .A1 (MultB_3), .A2 (nx1078), .B0 (
          nx954), .B1 (nx1080)) ;
    xnor2 ix1245 (.Y (nx1244), .A0 (nx1527), .A1 (nx1242)) ;
    nand02 ix1528 (.Y (nx1527), .A0 (MultA_11), .A1 (MultB_4)) ;
    xnor2 ix1243 (.Y (nx1242), .A0 (nx1531), .A1 (nx1240)) ;
    aoi32 ix1532 (.Y (nx1531), .A0 (MultA_10), .A1 (MultB_4), .A2 (nx1074), .B0 (
          nx962), .B1 (nx1076)) ;
    xnor2 ix1241 (.Y (nx1240), .A0 (nx1537), .A1 (nx1238)) ;
    nand02 ix1538 (.Y (nx1537), .A0 (MultA_10), .A1 (MultB_5)) ;
    xnor2 ix1239 (.Y (nx1238), .A0 (nx1541), .A1 (nx1236)) ;
    aoi32 ix1542 (.Y (nx1541), .A0 (MultA_9), .A1 (MultB_5), .A2 (nx1070), .B0 (
          nx970), .B1 (nx1072)) ;
    xnor2 ix1237 (.Y (nx1236), .A0 (nx1547), .A1 (nx1234)) ;
    nand02 ix1548 (.Y (nx1547), .A0 (MultA_9), .A1 (MultB_6)) ;
    xnor2 ix1235 (.Y (nx1234), .A0 (nx1551), .A1 (nx1232)) ;
    aoi32 ix1552 (.Y (nx1551), .A0 (MultA_8), .A1 (MultB_6), .A2 (nx1066), .B0 (
          nx978), .B1 (nx1068)) ;
    xnor2 ix1233 (.Y (nx1232), .A0 (nx1557), .A1 (nx1230)) ;
    nand02 ix1558 (.Y (nx1557), .A0 (MultA_8), .A1 (MultB_7)) ;
    xnor2 ix1231 (.Y (nx1230), .A0 (nx1561), .A1 (nx1228)) ;
    aoi32 ix1562 (.Y (nx1561), .A0 (MultA_7), .A1 (MultB_7), .A2 (nx1062), .B0 (
          nx986), .B1 (nx1064)) ;
    xnor2 ix1229 (.Y (nx1228), .A0 (nx1567), .A1 (nx1226)) ;
    nand02 ix1568 (.Y (nx1567), .A0 (MultA_7), .A1 (MultB_8)) ;
    xnor2 ix1227 (.Y (nx1226), .A0 (nx1571), .A1 (nx1224)) ;
    aoi32 ix1572 (.Y (nx1571), .A0 (MultA_6), .A1 (MultB_8), .A2 (nx1058), .B0 (
          nx994), .B1 (nx1060)) ;
    xnor2 ix1225 (.Y (nx1224), .A0 (nx1577), .A1 (nx1222)) ;
    nand02 ix1578 (.Y (nx1577), .A0 (MultA_6), .A1 (MultB_9)) ;
    xnor2 ix1223 (.Y (nx1222), .A0 (nx1581), .A1 (nx1220)) ;
    aoi32 ix1582 (.Y (nx1581), .A0 (MultA_5), .A1 (MultB_9), .A2 (nx1054), .B0 (
          nx1002), .B1 (nx1056)) ;
    xnor2 ix1221 (.Y (nx1220), .A0 (nx1587), .A1 (nx1218)) ;
    nand02 ix1588 (.Y (nx1587), .A0 (MultA_5), .A1 (MultB_10)) ;
    xnor2 ix1219 (.Y (nx1218), .A0 (nx1591), .A1 (nx1216)) ;
    aoi32 ix1592 (.Y (nx1591), .A0 (MultA_4), .A1 (MultB_10), .A2 (nx1050), .B0 (
          nx1010), .B1 (nx1052)) ;
    xnor2 ix1217 (.Y (nx1216), .A0 (nx1597), .A1 (nx1214)) ;
    nand02 ix1598 (.Y (nx1597), .A0 (MultA_4), .A1 (MultB_11)) ;
    xnor2 ix1215 (.Y (nx1214), .A0 (nx1601), .A1 (nx1212)) ;
    aoi32 ix1602 (.Y (nx1601), .A0 (MultA_3), .A1 (MultB_11), .A2 (nx1046), .B0 (
          nx1018), .B1 (nx1048)) ;
    xnor2 ix1213 (.Y (nx1212), .A0 (nx1607), .A1 (nx1210)) ;
    nand02 ix1608 (.Y (nx1607), .A0 (MultA_3), .A1 (MultB_12)) ;
    xnor2 ix1211 (.Y (nx1210), .A0 (nx1611), .A1 (nx1208)) ;
    aoi32 ix1612 (.Y (nx1611), .A0 (MultA_2), .A1 (MultB_12), .A2 (nx1042), .B0 (
          nx1026), .B1 (nx1044)) ;
    xnor2 ix1209 (.Y (nx1208), .A0 (nx1617), .A1 (nx1206)) ;
    nand02 ix1618 (.Y (nx1617), .A0 (MultA_2), .A1 (MultB_13)) ;
    xnor2 ix1207 (.Y (nx1206), .A0 (nx1198), .A1 (nx1631)) ;
    oai32 ix1199 (.Y (nx1198), .A0 (nx607), .A1 (nx1623), .A2 (nx1493), .B0 (
          nx1625), .B1 (nx1489)) ;
    inv01 ix1624 (.Y (nx1623), .A (MultB_13)) ;
    xnor2 ix1632 (.Y (nx1631), .A0 (nx1633), .A1 (nx1635)) ;
    nand02 ix1634 (.Y (nx1633), .A0 (MultA_1), .A1 (MultB_14)) ;
    nand02 ix1636 (.Y (nx1635), .A0 (MultB_15), .A1 (MultA_0)) ;
    mux21 ix2803 (.Y (Product_14), .A0 (nx1639), .A1 (nx2796), .S0 (nx509)) ;
    nand02 ix1640 (.Y (nx1639), .A0 (MultA_14), .A1 (MultB_0)) ;
    mux21 ix2811 (.Y (Product_13), .A0 (nx1645), .A1 (nx2804), .S0 (nx513)) ;
    nand02 ix1646 (.Y (nx1645), .A0 (MultA_13), .A1 (MultB_0)) ;
    mux21 ix2819 (.Y (Product_12), .A0 (nx1651), .A1 (nx2812), .S0 (nx517)) ;
    nand02 ix1652 (.Y (nx1651), .A0 (MultA_12), .A1 (MultB_0)) ;
    mux21 ix2827 (.Y (Product_11), .A0 (nx1657), .A1 (nx2820), .S0 (nx521)) ;
    nand02 ix1658 (.Y (nx1657), .A0 (MultA_11), .A1 (MultB_0)) ;
    mux21 ix2835 (.Y (Product_10), .A0 (nx1663), .A1 (nx2828), .S0 (nx525)) ;
    nand02 ix1664 (.Y (nx1663), .A0 (MultA_10), .A1 (MultB_0)) ;
    mux21 ix2843 (.Y (Product_9), .A0 (nx1669), .A1 (nx2836), .S0 (nx529)) ;
    nand02 ix1670 (.Y (nx1669), .A0 (MultA_9), .A1 (MultB_0)) ;
    mux21 ix2851 (.Y (Product_8), .A0 (nx1675), .A1 (nx2844), .S0 (nx533)) ;
    nand02 ix1676 (.Y (nx1675), .A0 (MultA_8), .A1 (MultB_0)) ;
    mux21 ix2859 (.Y (Product_7), .A0 (nx1681), .A1 (nx2852), .S0 (nx537)) ;
    nand02 ix1682 (.Y (nx1681), .A0 (MultA_7), .A1 (MultB_0)) ;
    mux21 ix2867 (.Y (Product_6), .A0 (nx1687), .A1 (nx2860), .S0 (nx541)) ;
    nand02 ix1688 (.Y (nx1687), .A0 (MultA_6), .A1 (MultB_0)) ;
    aoi21 ix2875 (.Y (Product_5), .A0 (nx1693), .A1 (nx545), .B0 (nx122)) ;
    nand02 ix1694 (.Y (nx1693), .A0 (MultA_5), .A1 (MultB_0)) ;
    aoi21 ix2883 (.Y (Product_4), .A0 (nx1697), .A1 (nx549), .B0 (nx74)) ;
    nand02 ix1698 (.Y (nx1697), .A0 (MultA_4), .A1 (MultB_0)) ;
    aoi21 ix2891 (.Y (Product_3), .A0 (nx1701), .A1 (nx553), .B0 (nx38)) ;
    nand02 ix1702 (.Y (nx1701), .A0 (MultA_3), .A1 (MultB_0)) ;
    aoi21 ix2899 (.Y (Product_2), .A0 (nx1705), .A1 (nx557), .B0 (nx14)) ;
    nand02 ix1706 (.Y (nx1705), .A0 (MultA_2), .A1 (MultB_0)) ;
    nor02ii ix2909 (.Y (Product_1), .A0 (nx1709), .A1 (nx559)) ;
    aoi22 ix1710 (.Y (nx1709), .A0 (MultA_1), .A1 (MultB_0), .B0 (MultB_1), .B1 (
          MultA_0)) ;
    xnor2 ix2787 (.Y (Product_16), .A0 (nx1262), .A1 (nx1715)) ;
    xnor2 ix1716 (.Y (nx1715), .A0 (nx1717), .A1 (nx1719)) ;
    nand02 ix1718 (.Y (nx1717), .A0 (MultA_15), .A1 (MultB_1)) ;
    xnor2 ix1720 (.Y (nx1719), .A0 (nx1721), .A1 (nx1723)) ;
    aoi32 ix1722 (.Y (nx1721), .A0 (MultA_14), .A1 (MultB_1), .A2 (nx1254), .B0 (
          nx1094), .B1 (nx1256)) ;
    xnor2 ix1724 (.Y (nx1723), .A0 (nx1725), .A1 (nx1727)) ;
    nand02 ix1726 (.Y (nx1725), .A0 (MultA_14), .A1 (MultB_2)) ;
    xnor2 ix1728 (.Y (nx1727), .A0 (nx1729), .A1 (nx1733)) ;
    aoi32 ix1730 (.Y (nx1729), .A0 (MultA_13), .A1 (MultB_2), .A2 (nx1250), .B0 (
          nx1102), .B1 (nx1252)) ;
    xnor2 ix1734 (.Y (nx1733), .A0 (nx1735), .A1 (nx1737)) ;
    nand02 ix1736 (.Y (nx1735), .A0 (MultA_13), .A1 (MultB_3)) ;
    xnor2 ix1738 (.Y (nx1737), .A0 (nx1739), .A1 (nx1743)) ;
    aoi32 ix1740 (.Y (nx1739), .A0 (MultA_12), .A1 (MultB_3), .A2 (nx1246), .B0 (
          nx1110), .B1 (nx1248)) ;
    xnor2 ix1744 (.Y (nx1743), .A0 (nx1745), .A1 (nx1747)) ;
    nand02 ix1746 (.Y (nx1745), .A0 (MultA_12), .A1 (MultB_4)) ;
    xnor2 ix1748 (.Y (nx1747), .A0 (nx1749), .A1 (nx1753)) ;
    aoi32 ix1750 (.Y (nx1749), .A0 (MultA_11), .A1 (MultB_4), .A2 (nx1242), .B0 (
          nx1118), .B1 (nx1244)) ;
    xnor2 ix1754 (.Y (nx1753), .A0 (nx1755), .A1 (nx1757)) ;
    nand02 ix1756 (.Y (nx1755), .A0 (MultA_11), .A1 (MultB_5)) ;
    xnor2 ix1758 (.Y (nx1757), .A0 (nx1759), .A1 (nx1763)) ;
    aoi32 ix1760 (.Y (nx1759), .A0 (MultA_10), .A1 (MultB_5), .A2 (nx1238), .B0 (
          nx1126), .B1 (nx1240)) ;
    xnor2 ix1764 (.Y (nx1763), .A0 (nx1765), .A1 (nx1767)) ;
    nand02 ix1766 (.Y (nx1765), .A0 (MultA_10), .A1 (MultB_6)) ;
    xnor2 ix1768 (.Y (nx1767), .A0 (nx1769), .A1 (nx1773)) ;
    aoi32 ix1770 (.Y (nx1769), .A0 (MultA_9), .A1 (MultB_6), .A2 (nx1234), .B0 (
          nx1134), .B1 (nx1236)) ;
    xnor2 ix1774 (.Y (nx1773), .A0 (nx1775), .A1 (nx1777)) ;
    nand02 ix1776 (.Y (nx1775), .A0 (MultA_9), .A1 (MultB_7)) ;
    xnor2 ix1778 (.Y (nx1777), .A0 (nx1779), .A1 (nx1783)) ;
    aoi32 ix1780 (.Y (nx1779), .A0 (MultA_8), .A1 (MultB_7), .A2 (nx1230), .B0 (
          nx1142), .B1 (nx1232)) ;
    xnor2 ix1784 (.Y (nx1783), .A0 (nx1785), .A1 (nx1787)) ;
    nand02 ix1786 (.Y (nx1785), .A0 (MultA_8), .A1 (MultB_8)) ;
    xnor2 ix1788 (.Y (nx1787), .A0 (nx1789), .A1 (nx1793)) ;
    aoi32 ix1790 (.Y (nx1789), .A0 (MultA_7), .A1 (MultB_8), .A2 (nx1226), .B0 (
          nx1150), .B1 (nx1228)) ;
    xnor2 ix1794 (.Y (nx1793), .A0 (nx1795), .A1 (nx1797)) ;
    nand02 ix1796 (.Y (nx1795), .A0 (MultA_7), .A1 (MultB_9)) ;
    xnor2 ix1798 (.Y (nx1797), .A0 (nx1799), .A1 (nx1803)) ;
    aoi32 ix1800 (.Y (nx1799), .A0 (MultA_6), .A1 (MultB_9), .A2 (nx1222), .B0 (
          nx1158), .B1 (nx1224)) ;
    xnor2 ix1804 (.Y (nx1803), .A0 (nx1805), .A1 (nx1807)) ;
    nand02 ix1806 (.Y (nx1805), .A0 (MultA_6), .A1 (MultB_10)) ;
    xnor2 ix1808 (.Y (nx1807), .A0 (nx1809), .A1 (nx1813)) ;
    aoi32 ix1810 (.Y (nx1809), .A0 (MultA_5), .A1 (MultB_10), .A2 (nx1218), .B0 (
          nx1166), .B1 (nx1220)) ;
    xnor2 ix1814 (.Y (nx1813), .A0 (nx1815), .A1 (nx1817)) ;
    nand02 ix1816 (.Y (nx1815), .A0 (MultA_5), .A1 (MultB_11)) ;
    xnor2 ix1818 (.Y (nx1817), .A0 (nx1819), .A1 (nx1823)) ;
    aoi32 ix1820 (.Y (nx1819), .A0 (MultA_4), .A1 (MultB_11), .A2 (nx1214), .B0 (
          nx1174), .B1 (nx1216)) ;
    xnor2 ix1824 (.Y (nx1823), .A0 (nx1825), .A1 (nx1827)) ;
    nand02 ix1826 (.Y (nx1825), .A0 (MultA_4), .A1 (MultB_12)) ;
    xnor2 ix1828 (.Y (nx1827), .A0 (nx1829), .A1 (nx1833)) ;
    aoi32 ix1830 (.Y (nx1829), .A0 (MultA_3), .A1 (MultB_12), .A2 (nx1210), .B0 (
          nx1182), .B1 (nx1212)) ;
    xnor2 ix1834 (.Y (nx1833), .A0 (nx1835), .A1 (nx1837)) ;
    nand02 ix1836 (.Y (nx1835), .A0 (MultA_3), .A1 (MultB_13)) ;
    xnor2 ix1838 (.Y (nx1837), .A0 (nx1839), .A1 (nx1843)) ;
    aoi32 ix1840 (.Y (nx1839), .A0 (MultA_2), .A1 (MultB_13), .A2 (nx1206), .B0 (
          nx1190), .B1 (nx1208)) ;
    xnor2 ix1844 (.Y (nx1843), .A0 (nx1845), .A1 (nx1847)) ;
    nand02 ix1846 (.Y (nx1845), .A0 (MultA_2), .A1 (MultB_14)) ;
    mux21 ix1848 (.Y (nx1847), .A0 (nx1849), .A1 (nx1376), .S0 (nx1374)) ;
    nand02 ix1850 (.Y (nx1849), .A0 (MultA_1), .A1 (MultB_15)) ;
    inv01 ix1854 (.Y (nx1853), .A (MultB_15)) ;
    oai32 ix1375 (.Y (nx1374), .A0 (nx607), .A1 (nx1857), .A2 (nx1635), .B0 (
          nx1859), .B1 (nx1631)) ;
    inv01 ix1858 (.Y (nx1857), .A (MultB_14)) ;
    xor2 ix2785 (.Y (Product_17), .A0 (nx1446), .A1 (nx1606)) ;
    xnor2 ix1607 (.Y (nx1606), .A0 (nx1873), .A1 (nx1604)) ;
    nand02 ix1874 (.Y (nx1873), .A0 (MultA_15), .A1 (MultB_2)) ;
    xnor2 ix1605 (.Y (nx1604), .A0 (nx1454), .A1 (nx1879)) ;
    oai32 ix1455 (.Y (nx1454), .A0 (nx1495), .A1 (nx609), .A2 (nx1727), .B0 (
          nx1721), .B1 (nx1723)) ;
    xnor2 ix1880 (.Y (nx1879), .A0 (nx1881), .A1 (nx1883)) ;
    nand02 ix1882 (.Y (nx1881), .A0 (MultA_14), .A1 (MultB_3)) ;
    xnor2 ix1884 (.Y (nx1883), .A0 (nx1462), .A1 (nx1598)) ;
    oai32 ix1463 (.Y (nx1462), .A0 (nx1363), .A1 (nx653), .A2 (nx1737), .B0 (
          nx1729), .B1 (nx1733)) ;
    xnor2 ix1599 (.Y (nx1598), .A0 (nx1889), .A1 (nx1596)) ;
    nand02 ix1890 (.Y (nx1889), .A0 (MultA_13), .A1 (MultB_4)) ;
    xnor2 ix1597 (.Y (nx1596), .A0 (nx1470), .A1 (nx1895)) ;
    oai32 ix1471 (.Y (nx1470), .A0 (nx1241), .A1 (nx705), .A2 (nx1747), .B0 (
          nx1739), .B1 (nx1743)) ;
    xnor2 ix1896 (.Y (nx1895), .A0 (nx1897), .A1 (nx1899)) ;
    nand02 ix1898 (.Y (nx1897), .A0 (MultA_12), .A1 (MultB_5)) ;
    xnor2 ix1900 (.Y (nx1899), .A0 (nx1478), .A1 (nx1590)) ;
    oai32 ix1479 (.Y (nx1478), .A0 (nx1129), .A1 (nx767), .A2 (nx1757), .B0 (
          nx1749), .B1 (nx1753)) ;
    xnor2 ix1591 (.Y (nx1590), .A0 (nx1905), .A1 (nx1588)) ;
    nand02 ix1906 (.Y (nx1905), .A0 (MultA_11), .A1 (MultB_6)) ;
    xnor2 ix1589 (.Y (nx1588), .A0 (nx1486), .A1 (nx1911)) ;
    oai32 ix1487 (.Y (nx1486), .A0 (nx1027), .A1 (nx839), .A2 (nx1767), .B0 (
          nx1759), .B1 (nx1763)) ;
    xnor2 ix1912 (.Y (nx1911), .A0 (nx1913), .A1 (nx1915)) ;
    nand02 ix1914 (.Y (nx1913), .A0 (MultA_10), .A1 (MultB_7)) ;
    xnor2 ix1916 (.Y (nx1915), .A0 (nx1494), .A1 (nx1582)) ;
    oai32 ix1495 (.Y (nx1494), .A0 (nx935), .A1 (nx921), .A2 (nx1777), .B0 (
          nx1769), .B1 (nx1773)) ;
    xnor2 ix1583 (.Y (nx1582), .A0 (nx1921), .A1 (nx1580)) ;
    nand02 ix1922 (.Y (nx1921), .A0 (MultA_9), .A1 (MultB_8)) ;
    xnor2 ix1581 (.Y (nx1580), .A0 (nx1502), .A1 (nx1927)) ;
    oai32 ix1503 (.Y (nx1502), .A0 (nx853), .A1 (nx1013), .A2 (nx1787), .B0 (
          nx1779), .B1 (nx1783)) ;
    xnor2 ix1928 (.Y (nx1927), .A0 (nx1929), .A1 (nx1931)) ;
    nand02 ix1930 (.Y (nx1929), .A0 (MultA_8), .A1 (MultB_9)) ;
    xnor2 ix1932 (.Y (nx1931), .A0 (nx1510), .A1 (nx1574)) ;
    oai32 ix1511 (.Y (nx1510), .A0 (nx781), .A1 (nx1115), .A2 (nx1797), .B0 (
          nx1789), .B1 (nx1793)) ;
    xnor2 ix1575 (.Y (nx1574), .A0 (nx1937), .A1 (nx1572)) ;
    nand02 ix1938 (.Y (nx1937), .A0 (MultA_7), .A1 (MultB_10)) ;
    xnor2 ix1573 (.Y (nx1572), .A0 (nx1518), .A1 (nx1943)) ;
    oai32 ix1519 (.Y (nx1518), .A0 (nx719), .A1 (nx1227), .A2 (nx1807), .B0 (
          nx1799), .B1 (nx1803)) ;
    xnor2 ix1944 (.Y (nx1943), .A0 (nx1945), .A1 (nx1947)) ;
    nand02 ix1946 (.Y (nx1945), .A0 (MultA_6), .A1 (MultB_11)) ;
    xnor2 ix1948 (.Y (nx1947), .A0 (nx1526), .A1 (nx1566)) ;
    oai32 ix1527 (.Y (nx1526), .A0 (nx667), .A1 (nx1349), .A2 (nx1817), .B0 (
          nx1809), .B1 (nx1813)) ;
    xnor2 ix1567 (.Y (nx1566), .A0 (nx1953), .A1 (nx1564)) ;
    nand02 ix1954 (.Y (nx1953), .A0 (MultA_5), .A1 (MultB_12)) ;
    xnor2 ix1565 (.Y (nx1564), .A0 (nx1534), .A1 (nx1959)) ;
    oai32 ix1535 (.Y (nx1534), .A0 (nx625), .A1 (nx1481), .A2 (nx1827), .B0 (
          nx1819), .B1 (nx1823)) ;
    xnor2 ix1960 (.Y (nx1959), .A0 (nx1961), .A1 (nx1963)) ;
    nand02 ix1962 (.Y (nx1961), .A0 (MultA_4), .A1 (MultB_13)) ;
    xnor2 ix1964 (.Y (nx1963), .A0 (nx1542), .A1 (nx1558)) ;
    oai32 ix1543 (.Y (nx1542), .A0 (nx589), .A1 (nx1623), .A2 (nx1837), .B0 (
          nx1829), .B1 (nx1833)) ;
    xnor2 ix1559 (.Y (nx1558), .A0 (nx1969), .A1 (nx1556)) ;
    nand02 ix1970 (.Y (nx1969), .A0 (MultA_3), .A1 (MultB_14)) ;
    xnor2 ix1557 (.Y (nx1556), .A0 (nx1550), .A1 (nx1975)) ;
    oai32 ix1551 (.Y (nx1550), .A0 (nx571), .A1 (nx1857), .A2 (nx1847), .B0 (
          nx1839), .B1 (nx1843)) ;
    xnor2 ix1976 (.Y (nx1975), .A0 (nx1977), .A1 (nx1979)) ;
    nand02 ix1978 (.Y (nx1977), .A0 (MultA_2), .A1 (MultB_15)) ;
    nand03 ix1980 (.Y (nx1979), .A0 (nx1374), .A1 (MultA_1), .A2 (MultB_15)) ;
    xnor2 ix2783 (.Y (Product_18), .A0 (nx1983), .A1 (nx1766)) ;
    aoi32 ix1984 (.Y (nx1983), .A0 (MultA_15), .A1 (MultB_2), .A2 (nx1604), .B0 (
          nx1446), .B1 (nx1606)) ;
    xnor2 ix1767 (.Y (nx1766), .A0 (nx1987), .A1 (nx1764)) ;
    nand02 ix1988 (.Y (nx1987), .A0 (MultA_15), .A1 (MultB_3)) ;
    xnor2 ix1765 (.Y (nx1764), .A0 (nx1620), .A1 (nx1995)) ;
    oai32 ix1621 (.Y (nx1620), .A0 (nx1495), .A1 (nx653), .A2 (nx1883), .B0 (
          nx1993), .B1 (nx1879)) ;
    inv01 ix1994 (.Y (nx1993), .A (nx1454)) ;
    xnor2 ix1996 (.Y (nx1995), .A0 (nx1997), .A1 (nx1999)) ;
    nand02 ix1998 (.Y (nx1997), .A0 (MultA_14), .A1 (MultB_4)) ;
    xnor2 ix2000 (.Y (nx1999), .A0 (nx2001), .A1 (nx2003)) ;
    aoi32 ix2002 (.Y (nx2001), .A0 (MultA_13), .A1 (MultB_4), .A2 (nx1596), .B0 (
          nx1462), .B1 (nx1598)) ;
    xnor2 ix2004 (.Y (nx2003), .A0 (nx2005), .A1 (nx2007)) ;
    nand02 ix2006 (.Y (nx2005), .A0 (MultA_13), .A1 (MultB_5)) ;
    xnor2 ix2008 (.Y (nx2007), .A0 (nx1636), .A1 (nx1754)) ;
    oai32 ix1637 (.Y (nx1636), .A0 (nx1241), .A1 (nx767), .A2 (nx1899), .B0 (
          nx2011), .B1 (nx1895)) ;
    inv01 ix2012 (.Y (nx2011), .A (nx1470)) ;
    xnor2 ix1755 (.Y (nx1754), .A0 (nx2015), .A1 (nx1752)) ;
    nand02 ix2016 (.Y (nx2015), .A0 (MultA_12), .A1 (MultB_6)) ;
    xnor2 ix1753 (.Y (nx1752), .A0 (nx2019), .A1 (nx1750)) ;
    aoi32 ix2020 (.Y (nx2019), .A0 (MultA_11), .A1 (MultB_6), .A2 (nx1588), .B0 (
          nx1478), .B1 (nx1590)) ;
    xnor2 ix1751 (.Y (nx1750), .A0 (nx2023), .A1 (nx1748)) ;
    nand02 ix2024 (.Y (nx2023), .A0 (MultA_11), .A1 (MultB_7)) ;
    xnor2 ix1749 (.Y (nx1748), .A0 (nx1652), .A1 (nx2031)) ;
    oai32 ix1653 (.Y (nx1652), .A0 (nx1027), .A1 (nx921), .A2 (nx1915), .B0 (
          nx2029), .B1 (nx1911)) ;
    inv01 ix2030 (.Y (nx2029), .A (nx1486)) ;
    xnor2 ix2032 (.Y (nx2031), .A0 (nx2033), .A1 (nx2035)) ;
    nand02 ix2034 (.Y (nx2033), .A0 (MultA_10), .A1 (MultB_8)) ;
    xnor2 ix2036 (.Y (nx2035), .A0 (nx2037), .A1 (nx2039)) ;
    aoi32 ix2038 (.Y (nx2037), .A0 (MultA_9), .A1 (MultB_8), .A2 (nx1580), .B0 (
          nx1494), .B1 (nx1582)) ;
    xnor2 ix2040 (.Y (nx2039), .A0 (nx2041), .A1 (nx2043)) ;
    nand02 ix2042 (.Y (nx2041), .A0 (MultA_9), .A1 (MultB_9)) ;
    xnor2 ix2044 (.Y (nx2043), .A0 (nx1668), .A1 (nx1738)) ;
    oai32 ix1669 (.Y (nx1668), .A0 (nx853), .A1 (nx1115), .A2 (nx1931), .B0 (
          nx2047), .B1 (nx1927)) ;
    inv01 ix2048 (.Y (nx2047), .A (nx1502)) ;
    xnor2 ix1739 (.Y (nx1738), .A0 (nx2051), .A1 (nx1736)) ;
    nand02 ix2052 (.Y (nx2051), .A0 (MultA_8), .A1 (MultB_10)) ;
    xnor2 ix1737 (.Y (nx1736), .A0 (nx2055), .A1 (nx1734)) ;
    aoi32 ix2056 (.Y (nx2055), .A0 (MultA_7), .A1 (MultB_10), .A2 (nx1572), .B0 (
          nx1510), .B1 (nx1574)) ;
    xnor2 ix1735 (.Y (nx1734), .A0 (nx2059), .A1 (nx1732)) ;
    nand02 ix2060 (.Y (nx2059), .A0 (MultA_7), .A1 (MultB_11)) ;
    xnor2 ix1733 (.Y (nx1732), .A0 (nx1684), .A1 (nx2067)) ;
    oai32 ix1685 (.Y (nx1684), .A0 (nx719), .A1 (nx1349), .A2 (nx1947), .B0 (
          nx2065), .B1 (nx1943)) ;
    inv01 ix2066 (.Y (nx2065), .A (nx1518)) ;
    xnor2 ix2068 (.Y (nx2067), .A0 (nx2069), .A1 (nx2071)) ;
    nand02 ix2070 (.Y (nx2069), .A0 (MultA_6), .A1 (MultB_12)) ;
    xnor2 ix2072 (.Y (nx2071), .A0 (nx2073), .A1 (nx2075)) ;
    aoi32 ix2074 (.Y (nx2073), .A0 (MultA_5), .A1 (MultB_12), .A2 (nx1564), .B0 (
          nx1526), .B1 (nx1566)) ;
    xnor2 ix2076 (.Y (nx2075), .A0 (nx2077), .A1 (nx2079)) ;
    nand02 ix2078 (.Y (nx2077), .A0 (MultA_5), .A1 (MultB_13)) ;
    xnor2 ix2080 (.Y (nx2079), .A0 (nx1700), .A1 (nx1722)) ;
    oai32 ix1701 (.Y (nx1700), .A0 (nx625), .A1 (nx1623), .A2 (nx1963), .B0 (
          nx2083), .B1 (nx1959)) ;
    inv01 ix2084 (.Y (nx2083), .A (nx1534)) ;
    xnor2 ix1723 (.Y (nx1722), .A0 (nx2087), .A1 (nx1720)) ;
    nand02 ix2088 (.Y (nx2087), .A0 (MultA_4), .A1 (MultB_14)) ;
    xnor2 ix1721 (.Y (nx1720), .A0 (nx2091), .A1 (nx1718)) ;
    aoi32 ix2092 (.Y (nx2091), .A0 (MultA_3), .A1 (MultB_14), .A2 (nx1556), .B0 (
          nx1542), .B1 (nx1558)) ;
    xnor2 ix1719 (.Y (nx1718), .A0 (nx2095), .A1 (nx1716)) ;
    nand02 ix2096 (.Y (nx2095), .A0 (MultA_3), .A1 (MultB_15)) ;
    oai32 ix1717 (.Y (nx1716), .A0 (nx571), .A1 (nx1853), .A2 (nx1979), .B0 (
          nx2099), .B1 (nx1975)) ;
    inv01 ix2100 (.Y (nx2099), .A (nx1550)) ;
    xor2 ix2781 (.Y (Product_19), .A0 (nx2103), .A1 (nx2107)) ;
    aoi32 ix2104 (.Y (nx2103), .A0 (MultA_15), .A1 (MultB_3), .A2 (nx1764), .B0 (
          nx1612), .B1 (nx1766)) ;
    xnor2 ix2108 (.Y (nx2107), .A0 (nx2109), .A1 (nx2111)) ;
    nand02 ix2110 (.Y (nx2109), .A0 (MultA_15), .A1 (MultB_4)) ;
    xnor2 ix2112 (.Y (nx2111), .A0 (nx1780), .A1 (nx1910)) ;
    oai32 ix1781 (.Y (nx1780), .A0 (nx1495), .A1 (nx705), .A2 (nx1999), .B0 (
          nx2115), .B1 (nx1995)) ;
    xnor2 ix1911 (.Y (nx1910), .A0 (nx2123), .A1 (nx1908)) ;
    nand02 ix2124 (.Y (nx2123), .A0 (MultA_14), .A1 (MultB_5)) ;
    xnor2 ix1909 (.Y (nx1908), .A0 (nx1788), .A1 (nx2129)) ;
    oai32 ix1789 (.Y (nx1788), .A0 (nx1363), .A1 (nx767), .A2 (nx2007), .B0 (
          nx2001), .B1 (nx2003)) ;
    xnor2 ix2130 (.Y (nx2129), .A0 (nx2131), .A1 (nx2133)) ;
    nand02 ix2132 (.Y (nx2131), .A0 (MultA_13), .A1 (MultB_6)) ;
    xnor2 ix2134 (.Y (nx2133), .A0 (nx2135), .A1 (nx2137)) ;
    aoi32 ix2136 (.Y (nx2135), .A0 (MultA_12), .A1 (MultB_6), .A2 (nx1752), .B0 (
          nx1636), .B1 (nx1754)) ;
    xnor2 ix2138 (.Y (nx2137), .A0 (nx2139), .A1 (nx2141)) ;
    nand02 ix2140 (.Y (nx2139), .A0 (MultA_12), .A1 (MultB_7)) ;
    xnor2 ix2142 (.Y (nx2141), .A0 (nx2143), .A1 (nx2147)) ;
    aoi32 ix2144 (.Y (nx2143), .A0 (MultA_11), .A1 (MultB_7), .A2 (nx1748), .B0 (
          nx1644), .B1 (nx1750)) ;
    xnor2 ix2148 (.Y (nx2147), .A0 (nx2149), .A1 (nx2151)) ;
    nand02 ix2150 (.Y (nx2149), .A0 (MultA_11), .A1 (MultB_8)) ;
    xnor2 ix2152 (.Y (nx2151), .A0 (nx1812), .A1 (nx1894)) ;
    oai32 ix1813 (.Y (nx1812), .A0 (nx1027), .A1 (nx1013), .A2 (nx2035), .B0 (
          nx2155), .B1 (nx2031)) ;
    xnor2 ix1895 (.Y (nx1894), .A0 (nx2163), .A1 (nx1892)) ;
    nand02 ix2164 (.Y (nx2163), .A0 (MultA_10), .A1 (MultB_9)) ;
    xnor2 ix1893 (.Y (nx1892), .A0 (nx1820), .A1 (nx2169)) ;
    oai32 ix1821 (.Y (nx1820), .A0 (nx935), .A1 (nx1115), .A2 (nx2043), .B0 (
          nx2037), .B1 (nx2039)) ;
    xnor2 ix2170 (.Y (nx2169), .A0 (nx2171), .A1 (nx2173)) ;
    nand02 ix2172 (.Y (nx2171), .A0 (MultA_9), .A1 (MultB_10)) ;
    xnor2 ix2174 (.Y (nx2173), .A0 (nx2175), .A1 (nx2177)) ;
    aoi32 ix2176 (.Y (nx2175), .A0 (MultA_8), .A1 (MultB_10), .A2 (nx1736), .B0 (
          nx1668), .B1 (nx1738)) ;
    xnor2 ix2178 (.Y (nx2177), .A0 (nx2179), .A1 (nx2181)) ;
    nand02 ix2180 (.Y (nx2179), .A0 (MultA_8), .A1 (MultB_11)) ;
    xnor2 ix2182 (.Y (nx2181), .A0 (nx2183), .A1 (nx2187)) ;
    aoi32 ix2184 (.Y (nx2183), .A0 (MultA_7), .A1 (MultB_11), .A2 (nx1732), .B0 (
          nx1676), .B1 (nx1734)) ;
    xnor2 ix2188 (.Y (nx2187), .A0 (nx2189), .A1 (nx2191)) ;
    nand02 ix2190 (.Y (nx2189), .A0 (MultA_7), .A1 (MultB_12)) ;
    xnor2 ix2192 (.Y (nx2191), .A0 (nx1844), .A1 (nx1878)) ;
    oai32 ix1845 (.Y (nx1844), .A0 (nx719), .A1 (nx1481), .A2 (nx2071), .B0 (
          nx2195), .B1 (nx2067)) ;
    xnor2 ix1879 (.Y (nx1878), .A0 (nx2203), .A1 (nx1876)) ;
    nand02 ix2204 (.Y (nx2203), .A0 (MultA_6), .A1 (MultB_13)) ;
    xnor2 ix1877 (.Y (nx1876), .A0 (nx1852), .A1 (nx2209)) ;
    oai32 ix1853 (.Y (nx1852), .A0 (nx667), .A1 (nx1623), .A2 (nx2079), .B0 (
          nx2073), .B1 (nx2075)) ;
    xnor2 ix2210 (.Y (nx2209), .A0 (nx2211), .A1 (nx2213)) ;
    nand02 ix2212 (.Y (nx2211), .A0 (MultA_5), .A1 (MultB_14)) ;
    xnor2 ix2214 (.Y (nx2213), .A0 (nx2215), .A1 (nx2217)) ;
    aoi32 ix2216 (.Y (nx2215), .A0 (MultA_4), .A1 (MultB_14), .A2 (nx1720), .B0 (
          nx1700), .B1 (nx1722)) ;
    xnor2 ix2218 (.Y (nx2217), .A0 (nx2219), .A1 (nx2221)) ;
    nand02 ix2220 (.Y (nx2219), .A0 (MultA_4), .A1 (MultB_15)) ;
    aoi32 ix2222 (.Y (nx2221), .A0 (MultA_3), .A1 (MultB_15), .A2 (nx1716), .B0 (
          nx1708), .B1 (nx1718)) ;
    xnor2 ix2779 (.Y (Product_20), .A0 (nx1920), .A1 (nx2229)) ;
    oai32 ix1921 (.Y (nx1920), .A0 (nx501), .A1 (nx705), .A2 (nx2111), .B0 (
          nx2103), .B1 (nx2107)) ;
    xnor2 ix2230 (.Y (nx2229), .A0 (nx2231), .A1 (nx2233)) ;
    nand02 ix2232 (.Y (nx2231), .A0 (MultA_15), .A1 (MultB_5)) ;
    xnor2 ix2234 (.Y (nx2233), .A0 (nx2235), .A1 (nx2237)) ;
    aoi32 ix2236 (.Y (nx2235), .A0 (MultA_14), .A1 (MultB_5), .A2 (nx1908), .B0 (
          nx1780), .B1 (nx1910)) ;
    xnor2 ix2238 (.Y (nx2237), .A0 (nx2239), .A1 (nx2241)) ;
    nand02 ix2240 (.Y (nx2239), .A0 (MultA_14), .A1 (MultB_6)) ;
    xnor2 ix2242 (.Y (nx2241), .A0 (nx1936), .A1 (nx2042)) ;
    oai32 ix1937 (.Y (nx1936), .A0 (nx1363), .A1 (nx839), .A2 (nx2133), .B0 (
          nx2245), .B1 (nx2129)) ;
    inv01 ix2246 (.Y (nx2245), .A (nx1788)) ;
    xnor2 ix2043 (.Y (nx2042), .A0 (nx2249), .A1 (nx2040)) ;
    nand02 ix2250 (.Y (nx2249), .A0 (MultA_13), .A1 (MultB_7)) ;
    xnor2 ix2041 (.Y (nx2040), .A0 (nx1944), .A1 (nx2255)) ;
    oai32 ix1945 (.Y (nx1944), .A0 (nx1241), .A1 (nx921), .A2 (nx2141), .B0 (
          nx2135), .B1 (nx2137)) ;
    xnor2 ix2256 (.Y (nx2255), .A0 (nx2257), .A1 (nx2259)) ;
    nand02 ix2258 (.Y (nx2257), .A0 (MultA_12), .A1 (MultB_8)) ;
    xnor2 ix2260 (.Y (nx2259), .A0 (nx1952), .A1 (nx2034)) ;
    oai32 ix1953 (.Y (nx1952), .A0 (nx1129), .A1 (nx1013), .A2 (nx2151), .B0 (
          nx2143), .B1 (nx2147)) ;
    xnor2 ix2035 (.Y (nx2034), .A0 (nx2265), .A1 (nx2032)) ;
    nand02 ix2266 (.Y (nx2265), .A0 (MultA_11), .A1 (MultB_9)) ;
    xnor2 ix2033 (.Y (nx2032), .A0 (nx2269), .A1 (nx2030)) ;
    aoi32 ix2270 (.Y (nx2269), .A0 (MultA_10), .A1 (MultB_9), .A2 (nx1892), .B0 (
          nx1812), .B1 (nx1894)) ;
    xnor2 ix2031 (.Y (nx2030), .A0 (nx2273), .A1 (nx2028)) ;
    nand02 ix2274 (.Y (nx2273), .A0 (MultA_10), .A1 (MultB_10)) ;
    xnor2 ix2029 (.Y (nx2028), .A0 (nx1968), .A1 (nx2281)) ;
    oai32 ix1969 (.Y (nx1968), .A0 (nx935), .A1 (nx1227), .A2 (nx2173), .B0 (
          nx2279), .B1 (nx2169)) ;
    inv01 ix2280 (.Y (nx2279), .A (nx1820)) ;
    xnor2 ix2282 (.Y (nx2281), .A0 (nx2283), .A1 (nx2285)) ;
    nand02 ix2284 (.Y (nx2283), .A0 (MultA_9), .A1 (MultB_11)) ;
    xnor2 ix2286 (.Y (nx2285), .A0 (nx1976), .A1 (nx2022)) ;
    oai32 ix1977 (.Y (nx1976), .A0 (nx853), .A1 (nx1349), .A2 (nx2181), .B0 (
          nx2175), .B1 (nx2177)) ;
    xnor2 ix2023 (.Y (nx2022), .A0 (nx2291), .A1 (nx2020)) ;
    nand02 ix2292 (.Y (nx2291), .A0 (MultA_8), .A1 (MultB_12)) ;
    xnor2 ix2021 (.Y (nx2020), .A0 (nx1984), .A1 (nx2297)) ;
    oai32 ix1985 (.Y (nx1984), .A0 (nx781), .A1 (nx1481), .A2 (nx2191), .B0 (
          nx2183), .B1 (nx2187)) ;
    xnor2 ix2298 (.Y (nx2297), .A0 (nx2299), .A1 (nx2301)) ;
    nand02 ix2300 (.Y (nx2299), .A0 (MultA_7), .A1 (MultB_13)) ;
    xnor2 ix2302 (.Y (nx2301), .A0 (nx2303), .A1 (nx2305)) ;
    aoi32 ix2304 (.Y (nx2303), .A0 (MultA_6), .A1 (MultB_13), .A2 (nx1876), .B0 (
          nx1844), .B1 (nx1878)) ;
    xnor2 ix2306 (.Y (nx2305), .A0 (nx2307), .A1 (nx2309)) ;
    nand02 ix2308 (.Y (nx2307), .A0 (MultA_6), .A1 (MultB_14)) ;
    xnor2 ix2310 (.Y (nx2309), .A0 (nx2000), .A1 (nx2010)) ;
    oai32 ix2001 (.Y (nx2000), .A0 (nx667), .A1 (nx1857), .A2 (nx2213), .B0 (
          nx2313), .B1 (nx2209)) ;
    inv01 ix2314 (.Y (nx2313), .A (nx1852)) ;
    xnor2 ix2011 (.Y (nx2010), .A0 (nx2317), .A1 (nx2008)) ;
    nand02 ix2318 (.Y (nx2317), .A0 (MultA_5), .A1 (MultB_15)) ;
    oai32 ix2009 (.Y (nx2008), .A0 (nx625), .A1 (nx1853), .A2 (nx2221), .B0 (
          nx2215), .B1 (nx2217)) ;
    xor2 ix2777 (.Y (Product_21), .A0 (nx2056), .A1 (nx2174)) ;
    oai32 ix2057 (.Y (nx2056), .A0 (nx501), .A1 (nx767), .A2 (nx2233), .B0 (
          nx2325), .B1 (nx2229)) ;
    inv01 ix2326 (.Y (nx2325), .A (nx1920)) ;
    xnor2 ix2175 (.Y (nx2174), .A0 (nx2329), .A1 (nx2172)) ;
    nand02 ix2330 (.Y (nx2329), .A0 (MultA_15), .A1 (MultB_6)) ;
    xnor2 ix2173 (.Y (nx2172), .A0 (nx2064), .A1 (nx2335)) ;
    oai32 ix2065 (.Y (nx2064), .A0 (nx1495), .A1 (nx839), .A2 (nx2241), .B0 (
          nx2235), .B1 (nx2237)) ;
    xnor2 ix2336 (.Y (nx2335), .A0 (nx2337), .A1 (nx2339)) ;
    nand02 ix2338 (.Y (nx2337), .A0 (MultA_14), .A1 (MultB_7)) ;
    xnor2 ix2340 (.Y (nx2339), .A0 (nx2341), .A1 (nx2343)) ;
    aoi32 ix2342 (.Y (nx2341), .A0 (MultA_13), .A1 (MultB_7), .A2 (nx2040), .B0 (
          nx1936), .B1 (nx2042)) ;
    xnor2 ix2344 (.Y (nx2343), .A0 (nx2345), .A1 (nx2347)) ;
    nand02 ix2346 (.Y (nx2345), .A0 (MultA_13), .A1 (MultB_8)) ;
    xnor2 ix2348 (.Y (nx2347), .A0 (nx2080), .A1 (nx2162)) ;
    oai32 ix2081 (.Y (nx2080), .A0 (nx1241), .A1 (nx1013), .A2 (nx2259), .B0 (
          nx2351), .B1 (nx2255)) ;
    inv01 ix2352 (.Y (nx2351), .A (nx1944)) ;
    xnor2 ix2163 (.Y (nx2162), .A0 (nx2355), .A1 (nx2160)) ;
    nand02 ix2356 (.Y (nx2355), .A0 (MultA_12), .A1 (MultB_9)) ;
    xnor2 ix2161 (.Y (nx2160), .A0 (nx2359), .A1 (nx2158)) ;
    aoi32 ix2360 (.Y (nx2359), .A0 (MultA_11), .A1 (MultB_9), .A2 (nx2032), .B0 (
          nx1952), .B1 (nx2034)) ;
    xnor2 ix2159 (.Y (nx2158), .A0 (nx2363), .A1 (nx2156)) ;
    nand02 ix2364 (.Y (nx2363), .A0 (MultA_11), .A1 (MultB_10)) ;
    xnor2 ix2157 (.Y (nx2156), .A0 (nx2367), .A1 (nx2154)) ;
    aoi32 ix2368 (.Y (nx2367), .A0 (MultA_10), .A1 (MultB_10), .A2 (nx2028), .B0 (
          nx1960), .B1 (nx2030)) ;
    xnor2 ix2155 (.Y (nx2154), .A0 (nx2373), .A1 (nx2152)) ;
    nand02 ix2374 (.Y (nx2373), .A0 (MultA_10), .A1 (MultB_11)) ;
    xnor2 ix2153 (.Y (nx2152), .A0 (nx2104), .A1 (nx2385)) ;
    oai32 ix2105 (.Y (nx2104), .A0 (nx935), .A1 (nx1349), .A2 (nx2285), .B0 (
          nx2379), .B1 (nx2281)) ;
    xnor2 ix2386 (.Y (nx2385), .A0 (nx2387), .A1 (nx2389)) ;
    nand02 ix2388 (.Y (nx2387), .A0 (MultA_9), .A1 (MultB_12)) ;
    xnor2 ix2390 (.Y (nx2389), .A0 (nx2391), .A1 (nx2393)) ;
    aoi32 ix2392 (.Y (nx2391), .A0 (MultA_8), .A1 (MultB_12), .A2 (nx2020), .B0 (
          nx1976), .B1 (nx2022)) ;
    xnor2 ix2394 (.Y (nx2393), .A0 (nx2395), .A1 (nx2397)) ;
    nand02 ix2396 (.Y (nx2395), .A0 (MultA_8), .A1 (MultB_13)) ;
    xnor2 ix2398 (.Y (nx2397), .A0 (nx2120), .A1 (nx2142)) ;
    oai32 ix2121 (.Y (nx2120), .A0 (nx781), .A1 (nx1623), .A2 (nx2301), .B0 (
          nx2401), .B1 (nx2297)) ;
    inv01 ix2402 (.Y (nx2401), .A (nx1984)) ;
    xnor2 ix2143 (.Y (nx2142), .A0 (nx2405), .A1 (nx2140)) ;
    nand02 ix2406 (.Y (nx2405), .A0 (MultA_7), .A1 (MultB_14)) ;
    xnor2 ix2141 (.Y (nx2140), .A0 (nx2128), .A1 (nx2411)) ;
    oai32 ix2129 (.Y (nx2128), .A0 (nx719), .A1 (nx1857), .A2 (nx2309), .B0 (
          nx2303), .B1 (nx2305)) ;
    xnor2 ix2412 (.Y (nx2411), .A0 (nx2413), .A1 (nx2415)) ;
    nand02 ix2414 (.Y (nx2413), .A0 (MultA_6), .A1 (MultB_15)) ;
    aoi32 ix2416 (.Y (nx2415), .A0 (MultA_5), .A1 (MultB_15), .A2 (nx2008), .B0 (
          nx2000), .B1 (nx2010)) ;
    xnor2 ix2775 (.Y (Product_22), .A0 (nx2419), .A1 (nx2286)) ;
    aoi32 ix2420 (.Y (nx2419), .A0 (MultA_15), .A1 (MultB_6), .A2 (nx2172), .B0 (
          nx2056), .B1 (nx2174)) ;
    xnor2 ix2287 (.Y (nx2286), .A0 (nx2423), .A1 (nx2284)) ;
    nand02 ix2424 (.Y (nx2423), .A0 (MultA_15), .A1 (MultB_7)) ;
    xnor2 ix2285 (.Y (nx2284), .A0 (nx2188), .A1 (nx2431)) ;
    oai32 ix2189 (.Y (nx2188), .A0 (nx1495), .A1 (nx921), .A2 (nx2339), .B0 (
          nx2429), .B1 (nx2335)) ;
    inv01 ix2430 (.Y (nx2429), .A (nx2064)) ;
    xnor2 ix2432 (.Y (nx2431), .A0 (nx2433), .A1 (nx2435)) ;
    nand02 ix2434 (.Y (nx2433), .A0 (MultA_14), .A1 (MultB_8)) ;
    xnor2 ix2436 (.Y (nx2435), .A0 (nx2196), .A1 (nx2278)) ;
    oai32 ix2197 (.Y (nx2196), .A0 (nx1363), .A1 (nx1013), .A2 (nx2347), .B0 (
          nx2341), .B1 (nx2343)) ;
    xnor2 ix2279 (.Y (nx2278), .A0 (nx2441), .A1 (nx2276)) ;
    nand02 ix2442 (.Y (nx2441), .A0 (MultA_13), .A1 (MultB_9)) ;
    xnor2 ix2277 (.Y (nx2276), .A0 (nx2445), .A1 (nx2274)) ;
    aoi32 ix2446 (.Y (nx2445), .A0 (MultA_12), .A1 (MultB_9), .A2 (nx2160), .B0 (
          nx2080), .B1 (nx2162)) ;
    xnor2 ix2275 (.Y (nx2274), .A0 (nx2449), .A1 (nx2272)) ;
    nand02 ix2450 (.Y (nx2449), .A0 (MultA_12), .A1 (MultB_10)) ;
    xnor2 ix2273 (.Y (nx2272), .A0 (nx2453), .A1 (nx2270)) ;
    aoi32 ix2454 (.Y (nx2453), .A0 (MultA_11), .A1 (MultB_10), .A2 (nx2156), .B0 (
          nx2088), .B1 (nx2158)) ;
    xnor2 ix2271 (.Y (nx2270), .A0 (nx2459), .A1 (nx2268)) ;
    nand02 ix2460 (.Y (nx2459), .A0 (MultA_11), .A1 (MultB_11)) ;
    xnor2 ix2269 (.Y (nx2268), .A0 (nx2463), .A1 (nx2266)) ;
    aoi32 ix2464 (.Y (nx2463), .A0 (MultA_10), .A1 (MultB_11), .A2 (nx2152), .B0 (
          nx2096), .B1 (nx2154)) ;
    xnor2 ix2267 (.Y (nx2266), .A0 (nx2469), .A1 (nx2264)) ;
    nand02 ix2470 (.Y (nx2469), .A0 (MultA_10), .A1 (MultB_12)) ;
    xnor2 ix2265 (.Y (nx2264), .A0 (nx2228), .A1 (nx2481)) ;
    oai32 ix2229 (.Y (nx2228), .A0 (nx935), .A1 (nx1481), .A2 (nx2389), .B0 (
          nx2475), .B1 (nx2385)) ;
    xnor2 ix2482 (.Y (nx2481), .A0 (nx2483), .A1 (nx2485)) ;
    nand02 ix2484 (.Y (nx2483), .A0 (MultA_9), .A1 (MultB_13)) ;
    xnor2 ix2486 (.Y (nx2485), .A0 (nx2236), .A1 (nx2258)) ;
    oai32 ix2237 (.Y (nx2236), .A0 (nx853), .A1 (nx1623), .A2 (nx2397), .B0 (
          nx2391), .B1 (nx2393)) ;
    xnor2 ix2259 (.Y (nx2258), .A0 (nx2491), .A1 (nx2256)) ;
    nand02 ix2492 (.Y (nx2491), .A0 (MultA_8), .A1 (MultB_14)) ;
    xnor2 ix2257 (.Y (nx2256), .A0 (nx2495), .A1 (nx2254)) ;
    aoi32 ix2496 (.Y (nx2495), .A0 (MultA_7), .A1 (MultB_14), .A2 (nx2140), .B0 (
          nx2120), .B1 (nx2142)) ;
    xnor2 ix2255 (.Y (nx2254), .A0 (nx2499), .A1 (nx2252)) ;
    nand02 ix2500 (.Y (nx2499), .A0 (MultA_7), .A1 (MultB_15)) ;
    oai32 ix2253 (.Y (nx2252), .A0 (nx719), .A1 (nx1853), .A2 (nx2415), .B0 (
          nx2503), .B1 (nx2411)) ;
    inv01 ix2504 (.Y (nx2503), .A (nx2128)) ;
    xor2 ix2773 (.Y (Product_23), .A0 (nx2507), .A1 (nx2511)) ;
    aoi32 ix2508 (.Y (nx2507), .A0 (MultA_15), .A1 (MultB_7), .A2 (nx2284), .B0 (
          nx2180), .B1 (nx2286)) ;
    xnor2 ix2512 (.Y (nx2511), .A0 (nx2513), .A1 (nx2515)) ;
    nand02 ix2514 (.Y (nx2513), .A0 (MultA_15), .A1 (MultB_8)) ;
    xnor2 ix2516 (.Y (nx2515), .A0 (nx2300), .A1 (nx2382)) ;
    oai32 ix2301 (.Y (nx2300), .A0 (nx1495), .A1 (nx1013), .A2 (nx2435), .B0 (
          nx2519), .B1 (nx2431)) ;
    xnor2 ix2383 (.Y (nx2382), .A0 (nx2527), .A1 (nx2380)) ;
    nand02 ix2528 (.Y (nx2527), .A0 (MultA_14), .A1 (MultB_9)) ;
    xnor2 ix2381 (.Y (nx2380), .A0 (nx2531), .A1 (nx2378)) ;
    aoi32 ix2532 (.Y (nx2531), .A0 (MultA_13), .A1 (MultB_9), .A2 (nx2276), .B0 (
          nx2196), .B1 (nx2278)) ;
    xnor2 ix2379 (.Y (nx2378), .A0 (nx2535), .A1 (nx2376)) ;
    nand02 ix2536 (.Y (nx2535), .A0 (MultA_13), .A1 (MultB_10)) ;
    xnor2 ix2377 (.Y (nx2376), .A0 (nx2539), .A1 (nx2374)) ;
    aoi32 ix2540 (.Y (nx2539), .A0 (MultA_12), .A1 (MultB_10), .A2 (nx2272), .B0 (
          nx2204), .B1 (nx2274)) ;
    xnor2 ix2375 (.Y (nx2374), .A0 (nx2545), .A1 (nx2372)) ;
    nand02 ix2546 (.Y (nx2545), .A0 (MultA_12), .A1 (MultB_11)) ;
    xnor2 ix2373 (.Y (nx2372), .A0 (nx2549), .A1 (nx2370)) ;
    aoi32 ix2550 (.Y (nx2549), .A0 (MultA_11), .A1 (MultB_11), .A2 (nx2268), .B0 (
          nx2212), .B1 (nx2270)) ;
    xnor2 ix2371 (.Y (nx2370), .A0 (nx2555), .A1 (nx2368)) ;
    nand02 ix2556 (.Y (nx2555), .A0 (MultA_11), .A1 (MultB_12)) ;
    xnor2 ix2369 (.Y (nx2368), .A0 (nx2559), .A1 (nx2366)) ;
    aoi32 ix2560 (.Y (nx2559), .A0 (MultA_10), .A1 (MultB_12), .A2 (nx2264), .B0 (
          nx2220), .B1 (nx2266)) ;
    xnor2 ix2367 (.Y (nx2366), .A0 (nx2565), .A1 (nx2364)) ;
    nand02 ix2566 (.Y (nx2565), .A0 (MultA_10), .A1 (MultB_13)) ;
    xnor2 ix2365 (.Y (nx2364), .A0 (nx2340), .A1 (nx2577)) ;
    oai32 ix2341 (.Y (nx2340), .A0 (nx935), .A1 (nx1623), .A2 (nx2485), .B0 (
          nx2571), .B1 (nx2481)) ;
    xnor2 ix2578 (.Y (nx2577), .A0 (nx2579), .A1 (nx2581)) ;
    nand02 ix2580 (.Y (nx2579), .A0 (MultA_9), .A1 (MultB_14)) ;
    xnor2 ix2582 (.Y (nx2581), .A0 (nx2583), .A1 (nx2585)) ;
    aoi32 ix2584 (.Y (nx2583), .A0 (MultA_8), .A1 (MultB_14), .A2 (nx2256), .B0 (
          nx2236), .B1 (nx2258)) ;
    xnor2 ix2586 (.Y (nx2585), .A0 (nx2587), .A1 (nx2589)) ;
    nand02 ix2588 (.Y (nx2587), .A0 (MultA_8), .A1 (MultB_15)) ;
    aoi32 ix2590 (.Y (nx2589), .A0 (MultA_7), .A1 (MultB_15), .A2 (nx2252), .B0 (
          nx2244), .B1 (nx2254)) ;
    xnor2 ix2771 (.Y (Product_24), .A0 (nx2392), .A1 (nx2597)) ;
    oai32 ix2393 (.Y (nx2392), .A0 (nx501), .A1 (nx1013), .A2 (nx2515), .B0 (
          nx2507), .B1 (nx2511)) ;
    xnor2 ix2598 (.Y (nx2597), .A0 (nx2599), .A1 (nx2601)) ;
    nand02 ix2600 (.Y (nx2599), .A0 (MultA_15), .A1 (MultB_9)) ;
    xnor2 ix2602 (.Y (nx2601), .A0 (nx2603), .A1 (nx2605)) ;
    aoi32 ix2604 (.Y (nx2603), .A0 (MultA_14), .A1 (MultB_9), .A2 (nx2380), .B0 (
          nx2300), .B1 (nx2382)) ;
    xnor2 ix2606 (.Y (nx2605), .A0 (nx2607), .A1 (nx2609)) ;
    nand02 ix2608 (.Y (nx2607), .A0 (MultA_14), .A1 (MultB_10)) ;
    xnor2 ix2610 (.Y (nx2609), .A0 (nx2611), .A1 (nx2615)) ;
    aoi32 ix2612 (.Y (nx2611), .A0 (MultA_13), .A1 (MultB_10), .A2 (nx2376), .B0 (
          nx2308), .B1 (nx2378)) ;
    xnor2 ix2616 (.Y (nx2615), .A0 (nx2617), .A1 (nx2619)) ;
    nand02 ix2618 (.Y (nx2617), .A0 (MultA_13), .A1 (MultB_11)) ;
    xnor2 ix2620 (.Y (nx2619), .A0 (nx2621), .A1 (nx2625)) ;
    aoi32 ix2622 (.Y (nx2621), .A0 (MultA_12), .A1 (MultB_11), .A2 (nx2372), .B0 (
          nx2316), .B1 (nx2374)) ;
    xnor2 ix2626 (.Y (nx2625), .A0 (nx2627), .A1 (nx2629)) ;
    nand02 ix2628 (.Y (nx2627), .A0 (MultA_12), .A1 (MultB_12)) ;
    xnor2 ix2630 (.Y (nx2629), .A0 (nx2631), .A1 (nx2635)) ;
    aoi32 ix2632 (.Y (nx2631), .A0 (MultA_11), .A1 (MultB_12), .A2 (nx2368), .B0 (
          nx2324), .B1 (nx2370)) ;
    xnor2 ix2636 (.Y (nx2635), .A0 (nx2637), .A1 (nx2639)) ;
    nand02 ix2638 (.Y (nx2637), .A0 (MultA_11), .A1 (MultB_13)) ;
    xnor2 ix2640 (.Y (nx2639), .A0 (nx2641), .A1 (nx2645)) ;
    aoi32 ix2642 (.Y (nx2641), .A0 (MultA_10), .A1 (MultB_13), .A2 (nx2364), .B0 (
          nx2332), .B1 (nx2366)) ;
    xnor2 ix2646 (.Y (nx2645), .A0 (nx2647), .A1 (nx2649)) ;
    nand02 ix2648 (.Y (nx2647), .A0 (MultA_10), .A1 (MultB_14)) ;
    xnor2 ix2650 (.Y (nx2649), .A0 (nx2440), .A1 (nx2450)) ;
    oai32 ix2441 (.Y (nx2440), .A0 (nx935), .A1 (nx1857), .A2 (nx2581), .B0 (
          nx2653), .B1 (nx2577)) ;
    xnor2 ix2451 (.Y (nx2450), .A0 (nx2661), .A1 (nx2448)) ;
    nand02 ix2662 (.Y (nx2661), .A0 (MultA_9), .A1 (MultB_15)) ;
    oai32 ix2449 (.Y (nx2448), .A0 (nx853), .A1 (nx1853), .A2 (nx2589), .B0 (
          nx2583), .B1 (nx2585)) ;
    xor2 ix2769 (.Y (Product_25), .A0 (nx2480), .A1 (nx2550)) ;
    oai32 ix2481 (.Y (nx2480), .A0 (nx501), .A1 (nx1115), .A2 (nx2601), .B0 (
          nx2669), .B1 (nx2597)) ;
    inv01 ix2670 (.Y (nx2669), .A (nx2392)) ;
    xnor2 ix2551 (.Y (nx2550), .A0 (nx2673), .A1 (nx2548)) ;
    nand02 ix2674 (.Y (nx2673), .A0 (MultA_15), .A1 (MultB_10)) ;
    xnor2 ix2549 (.Y (nx2548), .A0 (nx2488), .A1 (nx2679)) ;
    oai32 ix2489 (.Y (nx2488), .A0 (nx1495), .A1 (nx1227), .A2 (nx2609), .B0 (
          nx2603), .B1 (nx2605)) ;
    xnor2 ix2680 (.Y (nx2679), .A0 (nx2681), .A1 (nx2683)) ;
    nand02 ix2682 (.Y (nx2681), .A0 (MultA_14), .A1 (MultB_11)) ;
    xnor2 ix2684 (.Y (nx2683), .A0 (nx2496), .A1 (nx2542)) ;
    oai32 ix2497 (.Y (nx2496), .A0 (nx1363), .A1 (nx1349), .A2 (nx2619), .B0 (
          nx2611), .B1 (nx2615)) ;
    xnor2 ix2543 (.Y (nx2542), .A0 (nx2689), .A1 (nx2540)) ;
    nand02 ix2690 (.Y (nx2689), .A0 (MultA_13), .A1 (MultB_12)) ;
    xnor2 ix2541 (.Y (nx2540), .A0 (nx2504), .A1 (nx2695)) ;
    oai32 ix2505 (.Y (nx2504), .A0 (nx1241), .A1 (nx1481), .A2 (nx2629), .B0 (
          nx2621), .B1 (nx2625)) ;
    xnor2 ix2696 (.Y (nx2695), .A0 (nx2697), .A1 (nx2699)) ;
    nand02 ix2698 (.Y (nx2697), .A0 (MultA_12), .A1 (MultB_13)) ;
    xnor2 ix2700 (.Y (nx2699), .A0 (nx2512), .A1 (nx2534)) ;
    oai32 ix2513 (.Y (nx2512), .A0 (nx1129), .A1 (nx1623), .A2 (nx2639), .B0 (
          nx2631), .B1 (nx2635)) ;
    xnor2 ix2535 (.Y (nx2534), .A0 (nx2705), .A1 (nx2532)) ;
    nand02 ix2706 (.Y (nx2705), .A0 (MultA_11), .A1 (MultB_14)) ;
    xnor2 ix2533 (.Y (nx2532), .A0 (nx2520), .A1 (nx2711)) ;
    oai32 ix2521 (.Y (nx2520), .A0 (nx1027), .A1 (nx1857), .A2 (nx2649), .B0 (
          nx2641), .B1 (nx2645)) ;
    xnor2 ix2712 (.Y (nx2711), .A0 (nx2713), .A1 (nx2715)) ;
    nand02 ix2714 (.Y (nx2713), .A0 (MultA_10), .A1 (MultB_15)) ;
    aoi32 ix2716 (.Y (nx2715), .A0 (MultA_9), .A1 (MultB_15), .A2 (nx2448), .B0 (
          nx2440), .B1 (nx2450)) ;
    xnor2 ix2767 (.Y (Product_26), .A0 (nx2719), .A1 (nx2614)) ;
    aoi32 ix2720 (.Y (nx2719), .A0 (MultA_15), .A1 (MultB_10), .A2 (nx2548), .B0 (
          nx2480), .B1 (nx2550)) ;
    xnor2 ix2615 (.Y (nx2614), .A0 (nx2723), .A1 (nx2612)) ;
    nand02 ix2724 (.Y (nx2723), .A0 (MultA_15), .A1 (MultB_11)) ;
    xnor2 ix2613 (.Y (nx2612), .A0 (nx2564), .A1 (nx2731)) ;
    oai32 ix2565 (.Y (nx2564), .A0 (nx1495), .A1 (nx1349), .A2 (nx2683), .B0 (
          nx2729), .B1 (nx2679)) ;
    inv01 ix2730 (.Y (nx2729), .A (nx2488)) ;
    xnor2 ix2732 (.Y (nx2731), .A0 (nx2733), .A1 (nx2735)) ;
    nand02 ix2734 (.Y (nx2733), .A0 (MultA_14), .A1 (MultB_12)) ;
    xnor2 ix2736 (.Y (nx2735), .A0 (nx2737), .A1 (nx2739)) ;
    aoi32 ix2738 (.Y (nx2737), .A0 (MultA_13), .A1 (MultB_12), .A2 (nx2540), .B0 (
          nx2496), .B1 (nx2542)) ;
    xnor2 ix2740 (.Y (nx2739), .A0 (nx2741), .A1 (nx2743)) ;
    nand02 ix2742 (.Y (nx2741), .A0 (MultA_13), .A1 (MultB_13)) ;
    xnor2 ix2744 (.Y (nx2743), .A0 (nx2580), .A1 (nx2602)) ;
    oai32 ix2581 (.Y (nx2580), .A0 (nx1241), .A1 (nx1623), .A2 (nx2699), .B0 (
          nx2747), .B1 (nx2695)) ;
    inv01 ix2748 (.Y (nx2747), .A (nx2504)) ;
    xnor2 ix2603 (.Y (nx2602), .A0 (nx2751), .A1 (nx2600)) ;
    nand02 ix2752 (.Y (nx2751), .A0 (MultA_12), .A1 (MultB_14)) ;
    xnor2 ix2601 (.Y (nx2600), .A0 (nx2755), .A1 (nx2598)) ;
    aoi32 ix2756 (.Y (nx2755), .A0 (MultA_11), .A1 (MultB_14), .A2 (nx2532), .B0 (
          nx2512), .B1 (nx2534)) ;
    xnor2 ix2599 (.Y (nx2598), .A0 (nx2759), .A1 (nx2596)) ;
    nand02 ix2760 (.Y (nx2759), .A0 (MultA_11), .A1 (MultB_15)) ;
    oai32 ix2597 (.Y (nx2596), .A0 (nx1027), .A1 (nx1853), .A2 (nx2715), .B0 (
          nx2763), .B1 (nx2711)) ;
    inv01 ix2764 (.Y (nx2763), .A (nx2520)) ;
    xor2 ix2765 (.Y (Product_27), .A0 (nx2767), .A1 (nx2771)) ;
    aoi32 ix2768 (.Y (nx2767), .A0 (MultA_15), .A1 (MultB_11), .A2 (nx2612), .B0 (
          nx2556), .B1 (nx2614)) ;
    xnor2 ix2772 (.Y (nx2771), .A0 (nx2773), .A1 (nx2775)) ;
    nand02 ix2774 (.Y (nx2773), .A0 (MultA_15), .A1 (MultB_12)) ;
    xnor2 ix2776 (.Y (nx2775), .A0 (nx2628), .A1 (nx2662)) ;
    oai32 ix2629 (.Y (nx2628), .A0 (nx1495), .A1 (nx1481), .A2 (nx2735), .B0 (
          nx2779), .B1 (nx2731)) ;
    xnor2 ix2663 (.Y (nx2662), .A0 (nx2787), .A1 (nx2660)) ;
    nand02 ix2788 (.Y (nx2787), .A0 (MultA_14), .A1 (MultB_13)) ;
    xnor2 ix2661 (.Y (nx2660), .A0 (nx2636), .A1 (nx2793)) ;
    oai32 ix2637 (.Y (nx2636), .A0 (nx1363), .A1 (nx1623), .A2 (nx2743), .B0 (
          nx2737), .B1 (nx2739)) ;
    xnor2 ix2794 (.Y (nx2793), .A0 (nx2795), .A1 (nx2797)) ;
    nand02 ix2796 (.Y (nx2795), .A0 (MultA_13), .A1 (MultB_14)) ;
    xnor2 ix2798 (.Y (nx2797), .A0 (nx2799), .A1 (nx2801)) ;
    aoi32 ix2800 (.Y (nx2799), .A0 (MultA_12), .A1 (MultB_14), .A2 (nx2600), .B0 (
          nx2580), .B1 (nx2602)) ;
    xnor2 ix2802 (.Y (nx2801), .A0 (nx2803), .A1 (nx2805)) ;
    nand02 ix2804 (.Y (nx2803), .A0 (MultA_12), .A1 (MultB_15)) ;
    aoi32 ix2806 (.Y (nx2805), .A0 (MultA_11), .A1 (MultB_15), .A2 (nx2596), .B0 (
          nx2588), .B1 (nx2598)) ;
    xnor2 ix2763 (.Y (Product_28), .A0 (nx2672), .A1 (nx2813)) ;
    oai32 ix2673 (.Y (nx2672), .A0 (nx501), .A1 (nx1481), .A2 (nx2775), .B0 (
          nx2767), .B1 (nx2771)) ;
    xnor2 ix2814 (.Y (nx2813), .A0 (nx2815), .A1 (nx2817)) ;
    nand02 ix2816 (.Y (nx2815), .A0 (MultA_15), .A1 (MultB_13)) ;
    xnor2 ix2818 (.Y (nx2817), .A0 (nx2819), .A1 (nx2821)) ;
    aoi32 ix2820 (.Y (nx2819), .A0 (MultA_14), .A1 (MultB_13), .A2 (nx2660), .B0 (
          nx2628), .B1 (nx2662)) ;
    xnor2 ix2822 (.Y (nx2821), .A0 (nx2823), .A1 (nx2825)) ;
    nand02 ix2824 (.Y (nx2823), .A0 (MultA_14), .A1 (MultB_14)) ;
    xnor2 ix2826 (.Y (nx2825), .A0 (nx2688), .A1 (nx2698)) ;
    oai32 ix2689 (.Y (nx2688), .A0 (nx1363), .A1 (nx1857), .A2 (nx2797), .B0 (
          nx2829), .B1 (nx2793)) ;
    inv01 ix2830 (.Y (nx2829), .A (nx2636)) ;
    xnor2 ix2699 (.Y (nx2698), .A0 (nx2833), .A1 (nx2696)) ;
    nand02 ix2834 (.Y (nx2833), .A0 (MultA_13), .A1 (MultB_15)) ;
    oai32 ix2697 (.Y (nx2696), .A0 (nx1241), .A1 (nx1853), .A2 (nx2805), .B0 (
          nx2799), .B1 (nx2801)) ;
    xor2 ix2761 (.Y (Product_29), .A0 (nx2712), .A1 (nx2734)) ;
    oai32 ix2713 (.Y (nx2712), .A0 (nx501), .A1 (nx1623), .A2 (nx2817), .B0 (
          nx2841), .B1 (nx2813)) ;
    inv01 ix2842 (.Y (nx2841), .A (nx2672)) ;
    xnor2 ix2735 (.Y (nx2734), .A0 (nx2845), .A1 (nx2732)) ;
    nand02 ix2846 (.Y (nx2845), .A0 (MultA_15), .A1 (MultB_14)) ;
    xnor2 ix2733 (.Y (nx2732), .A0 (nx2720), .A1 (nx2851)) ;
    oai32 ix2721 (.Y (nx2720), .A0 (nx1495), .A1 (nx1857), .A2 (nx2825), .B0 (
          nx2819), .B1 (nx2821)) ;
    xnor2 ix2852 (.Y (nx2851), .A0 (nx2853), .A1 (nx2855)) ;
    nand02 ix2854 (.Y (nx2853), .A0 (MultA_14), .A1 (MultB_15)) ;
    aoi32 ix2856 (.Y (nx2855), .A0 (MultA_13), .A1 (MultB_15), .A2 (nx2696), .B0 (
          nx2688), .B1 (nx2698)) ;
    xnor2 ix2759 (.Y (Product_30), .A0 (nx2859), .A1 (nx2750)) ;
    aoi32 ix2860 (.Y (nx2859), .A0 (MultA_15), .A1 (MultB_14), .A2 (nx2732), .B0 (
          nx2712), .B1 (nx2734)) ;
    xnor2 ix2751 (.Y (nx2750), .A0 (nx2863), .A1 (nx2748)) ;
    nand02 ix2864 (.Y (nx2863), .A0 (MultA_15), .A1 (MultB_15)) ;
    oai32 ix2749 (.Y (nx2748), .A0 (nx1495), .A1 (nx1853), .A2 (nx2855), .B0 (
          nx2867), .B1 (nx2851)) ;
    inv01 ix2868 (.Y (nx2867), .A (nx2720)) ;
    ao32 ix2757 (.Y (Product_31), .A0 (MultA_15), .A1 (MultB_15), .A2 (nx2748), 
         .B0 (nx2740), .B1 (nx2750)) ;
    inv01 ix2741 (.Y (nx2740), .A (nx2859)) ;
    inv01 ix2589 (.Y (nx2588), .A (nx2755)) ;
    inv01 ix2780 (.Y (nx2779), .A (nx2564)) ;
    inv01 ix2557 (.Y (nx2556), .A (nx2719)) ;
    inv01 ix2654 (.Y (nx2653), .A (nx2340)) ;
    inv01 ix2333 (.Y (nx2332), .A (nx2559)) ;
    inv01 ix2325 (.Y (nx2324), .A (nx2549)) ;
    inv01 ix2317 (.Y (nx2316), .A (nx2539)) ;
    inv01 ix2309 (.Y (nx2308), .A (nx2531)) ;
    inv01 ix2245 (.Y (nx2244), .A (nx2495)) ;
    inv01 ix2572 (.Y (nx2571), .A (nx2228)) ;
    inv01 ix2221 (.Y (nx2220), .A (nx2463)) ;
    inv01 ix2213 (.Y (nx2212), .A (nx2453)) ;
    inv01 ix2205 (.Y (nx2204), .A (nx2445)) ;
    inv01 ix2520 (.Y (nx2519), .A (nx2188)) ;
    inv01 ix2181 (.Y (nx2180), .A (nx2419)) ;
    inv01 ix2476 (.Y (nx2475), .A (nx2104)) ;
    inv01 ix2097 (.Y (nx2096), .A (nx2367)) ;
    inv01 ix2089 (.Y (nx2088), .A (nx2359)) ;
    inv01 ix2380 (.Y (nx2379), .A (nx1968)) ;
    inv01 ix1961 (.Y (nx1960), .A (nx2269)) ;
    inv01 ix1709 (.Y (nx1708), .A (nx2091)) ;
    inv01 ix2196 (.Y (nx2195), .A (nx1684)) ;
    inv01 ix1677 (.Y (nx1676), .A (nx2055)) ;
    inv01 ix2156 (.Y (nx2155), .A (nx1652)) ;
    inv01 ix1645 (.Y (nx1644), .A (nx2019)) ;
    inv01 ix2116 (.Y (nx2115), .A (nx1620)) ;
    inv01 ix1613 (.Y (nx1612), .A (nx1983)) ;
    inv01 ix1860 (.Y (nx1859), .A (nx1198)) ;
    inv01 ix1191 (.Y (nx1190), .A (nx1611)) ;
    inv01 ix1183 (.Y (nx1182), .A (nx1601)) ;
    inv01 ix1175 (.Y (nx1174), .A (nx1591)) ;
    inv01 ix1167 (.Y (nx1166), .A (nx1581)) ;
    inv01 ix1159 (.Y (nx1158), .A (nx1571)) ;
    inv01 ix1151 (.Y (nx1150), .A (nx1561)) ;
    inv01 ix1143 (.Y (nx1142), .A (nx1551)) ;
    inv01 ix1135 (.Y (nx1134), .A (nx1541)) ;
    inv01 ix1127 (.Y (nx1126), .A (nx1531)) ;
    inv01 ix1119 (.Y (nx1118), .A (nx1521)) ;
    inv01 ix1111 (.Y (nx1110), .A (nx1511)) ;
    inv01 ix1103 (.Y (nx1102), .A (nx1503)) ;
    inv01 ix1626 (.Y (nx1625), .A (nx1034)) ;
    inv01 ix1027 (.Y (nx1026), .A (nx1469)) ;
    inv01 ix1019 (.Y (nx1018), .A (nx1459)) ;
    inv01 ix1011 (.Y (nx1010), .A (nx1449)) ;
    inv01 ix1003 (.Y (nx1002), .A (nx1439)) ;
    inv01 ix995 (.Y (nx994), .A (nx1429)) ;
    inv01 ix987 (.Y (nx986), .A (nx1419)) ;
    inv01 ix979 (.Y (nx978), .A (nx1409)) ;
    inv01 ix971 (.Y (nx970), .A (nx1399)) ;
    inv01 ix963 (.Y (nx962), .A (nx1389)) ;
    inv01 ix955 (.Y (nx954), .A (nx1379)) ;
    inv01 ix947 (.Y (nx946), .A (nx1371)) ;
    inv01 ix1484 (.Y (nx1483), .A (nx882)) ;
    inv01 ix875 (.Y (nx874), .A (nx1337)) ;
    inv01 ix867 (.Y (nx866), .A (nx1327)) ;
    inv01 ix859 (.Y (nx858), .A (nx1317)) ;
    inv01 ix851 (.Y (nx850), .A (nx1307)) ;
    inv01 ix843 (.Y (nx842), .A (nx1297)) ;
    inv01 ix835 (.Y (nx834), .A (nx1287)) ;
    inv01 ix827 (.Y (nx826), .A (nx1277)) ;
    inv01 ix819 (.Y (nx818), .A (nx1267)) ;
    inv01 ix811 (.Y (nx810), .A (nx1257)) ;
    inv01 ix803 (.Y (nx802), .A (nx1249)) ;
    inv01 ix1352 (.Y (nx1351), .A (nx742)) ;
    inv01 ix735 (.Y (nx734), .A (nx1215)) ;
    inv01 ix727 (.Y (nx726), .A (nx1205)) ;
    inv01 ix719 (.Y (nx718), .A (nx1195)) ;
    inv01 ix711 (.Y (nx710), .A (nx1185)) ;
    inv01 ix703 (.Y (nx702), .A (nx1175)) ;
    inv01 ix695 (.Y (nx694), .A (nx1165)) ;
    inv01 ix687 (.Y (nx686), .A (nx1155)) ;
    inv01 ix679 (.Y (nx678), .A (nx1145)) ;
    inv01 ix671 (.Y (nx670), .A (nx1137)) ;
    inv01 ix1230 (.Y (nx1229), .A (nx614)) ;
    inv01 ix607 (.Y (nx606), .A (nx1103)) ;
    inv01 ix599 (.Y (nx598), .A (nx1093)) ;
    inv01 ix591 (.Y (nx590), .A (nx1083)) ;
    inv01 ix583 (.Y (nx582), .A (nx1073)) ;
    inv01 ix575 (.Y (nx574), .A (nx1063)) ;
    inv01 ix567 (.Y (nx566), .A (nx1053)) ;
    inv01 ix559 (.Y (nx558), .A (nx1043)) ;
    inv01 ix551 (.Y (nx550), .A (nx1035)) ;
    inv01 ix1118 (.Y (nx1117), .A (nx498)) ;
    inv01 ix491 (.Y (nx490), .A (nx1001)) ;
    inv01 ix483 (.Y (nx482), .A (nx991)) ;
    inv01 ix475 (.Y (nx474), .A (nx981)) ;
    inv01 ix467 (.Y (nx466), .A (nx971)) ;
    inv01 ix459 (.Y (nx458), .A (nx961)) ;
    inv01 ix451 (.Y (nx450), .A (nx951)) ;
    inv01 ix443 (.Y (nx442), .A (nx943)) ;
    inv01 ix1016 (.Y (nx1015), .A (nx394)) ;
    inv01 ix387 (.Y (nx386), .A (nx909)) ;
    inv01 ix379 (.Y (nx378), .A (nx899)) ;
    inv01 ix371 (.Y (nx370), .A (nx889)) ;
    inv01 ix363 (.Y (nx362), .A (nx879)) ;
    inv01 ix355 (.Y (nx354), .A (nx869)) ;
    inv01 ix347 (.Y (nx346), .A (nx861)) ;
    inv01 ix924 (.Y (nx923), .A (nx302)) ;
    inv01 ix295 (.Y (nx294), .A (nx827)) ;
    inv01 ix287 (.Y (nx286), .A (nx817)) ;
    inv01 ix279 (.Y (nx278), .A (nx807)) ;
    inv01 ix271 (.Y (nx270), .A (nx797)) ;
    inv01 ix263 (.Y (nx262), .A (nx789)) ;
    inv01 ix842 (.Y (nx841), .A (nx222)) ;
    inv01 ix215 (.Y (nx214), .A (nx755)) ;
    inv01 ix207 (.Y (nx206), .A (nx745)) ;
    inv01 ix199 (.Y (nx198), .A (nx735)) ;
    inv01 ix191 (.Y (nx190), .A (nx727)) ;
    inv01 ix770 (.Y (nx769), .A (nx154)) ;
    inv01 ix147 (.Y (nx146), .A (nx693)) ;
    inv01 ix139 (.Y (nx138), .A (nx683)) ;
    inv01 ix131 (.Y (nx130), .A (nx675)) ;
    inv01 ix708 (.Y (nx707), .A (nx98)) ;
    inv01 ix91 (.Y (nx90), .A (nx641)) ;
    inv01 ix83 (.Y (nx82), .A (nx633)) ;
    inv01 ix656 (.Y (nx655), .A (nx54)) ;
    inv01 ix47 (.Y (nx46), .A (nx597)) ;
    inv01 ix612 (.Y (nx611), .A (nx22)) ;
    inv01 ix3 (.Y (Product_0), .A (nx581)) ;
    inv02 ix2877 (.Y (nx2878), .A (MultB_0)) ;
    and02 ix2789 (.Y (nx2788), .A0 (MultA_15), .A1 (MultB_0)) ;
    and02 ix2797 (.Y (nx2796), .A0 (MultA_14), .A1 (MultB_0)) ;
    and02 ix2805 (.Y (nx2804), .A0 (MultA_13), .A1 (MultB_0)) ;
    and02 ix2813 (.Y (nx2812), .A0 (MultA_12), .A1 (MultB_0)) ;
    and02 ix2821 (.Y (nx2820), .A0 (MultA_11), .A1 (MultB_0)) ;
    and02 ix2829 (.Y (nx2828), .A0 (MultA_10), .A1 (MultB_0)) ;
    and02 ix2837 (.Y (nx2836), .A0 (MultA_9), .A1 (MultB_0)) ;
    and02 ix2845 (.Y (nx2844), .A0 (MultA_8), .A1 (MultB_0)) ;
    and02 ix2853 (.Y (nx2852), .A0 (MultA_7), .A1 (MultB_0)) ;
    and02 ix2861 (.Y (nx2860), .A0 (MultA_6), .A1 (MultB_0)) ;
    and03 ix1263 (.Y (nx1262), .A0 (nx2886), .A1 (MultA_15), .A2 (MultB_0)) ;
    inv01 ix2885 (.Y (nx2886), .A (nx505)) ;
    and02 ix1377 (.Y (nx1376), .A0 (MultA_1), .A1 (MultB_15)) ;
    ao32 ix1447 (.Y (nx1446), .A0 (MultA_15), .A1 (MultB_1), .A2 (nx2888), .B0 (
         nx1262), .B1 (nx2890)) ;
    inv01 ix2887 (.Y (nx2888), .A (nx1719)) ;
    inv01 ix2889 (.Y (nx2890), .A (nx1715)) ;
endmodule


module full_adder ( A, B, Cin, Sum, Cout ) ;

    input A ;
    input B ;
    input Cin ;
    output Sum ;
    output Cout ;




endmodule


module nBitRegister_32 ( nBitIn, WE, Reset, clk, Y ) ;

    input [31:0]nBitIn ;
    input WE ;
    input Reset ;
    input clk ;
    output [31:0]Y ;




endmodule


module nBitRegister_16 ( nBitIn, WE, Reset, clk, Y ) ;

    input [15:0]nBitIn ;
    input WE ;
    input Reset ;
    input clk ;
    output [15:0]Y ;




endmodule

