
-- 
-- Definition of  ProjectWrapper
-- 
--      Mon Nov 25 19:21:25 2019
--      
--      LeonardoSpectrum Level 3, 2008b.3
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity ProjectWrapper is
   port (
      A : IN std_logic_vector (15 DOWNTO 0) ;
      B : IN std_logic_vector (15 DOWNTO 0) ;
      clk : IN std_logic ;
      WE : IN std_logic ;
      reset : IN std_logic ;
      StartTest : IN std_logic ;
      RegOut : OUT std_logic_vector (31 DOWNTO 0) ;
      Pass : OUT std_logic ;
      Complete : OUT std_logic) ;
end ProjectWrapper ;

architecture Behavioral of ProjectWrapper is
   signal RegOut_dup0_31, RegOut_dup0_30, RegOut_dup0_29, RegOut_dup0_28, 
      RegOut_dup0_27, RegOut_dup0_26, RegOut_dup0_25, RegOut_dup0_24, 
      RegOut_dup0_23, RegOut_dup0_22, RegOut_dup0_21, RegOut_dup0_20, 
      RegOut_dup0_19, RegOut_dup0_18, RegOut_dup0_17, RegOut_dup0_16, 
      RegOut_dup0_15, RegOut_dup0_14, RegOut_dup0_13, RegOut_dup0_12, 
      RegOut_dup0_11, RegOut_dup0_10, RegOut_dup0_9, RegOut_dup0_8, 
      RegOut_dup0_7, RegOut_dup0_6, RegOut_dup0_5, RegOut_dup0_4, 
      RegOut_dup0_3, RegOut_dup0_2, RegOut_dup0_1, RegOut_dup0_0, Pass_dup0, 
      Complete_dup0, CounterOut_31, CounterOut_30, CounterOut_29, nx935, 
      CounterOut_28, CounterOut_27, nx939, CounterOut_26, CounterOut_25, 
      nx943, CounterOut_24, CounterOut_23, nx947, CounterOut_22, 
      CounterOut_21, nx951, CounterOut_20, CounterOut_19, nx955, 
      CounterOut_18, CounterOut_17, nx959, CounterOut_16, CounterOut_15, 
      nx963, CounterOut_14, CounterOut_13, nx965, CounterOut_12, 
      CounterOut_11, nx967, CounterOut_10, CounterOut_9, nx971, CounterOut_8, 
      CounterOut_7, nx975, CounterOut_6, CounterOut_5, nx979, CounterOut_4, 
      CounterOut_3, nx983, CounterOut_2, nx985, CounterOut_1, nx987, 
      CounterOut_0, nx30, nx44, nx58, nx72, nx86, nx100, nx114, nx128, nx142, 
      nx156, nx170, nx184, nx198, nx212, nx226, nx240, nx254, nx268, nx282, 
      nx296, nx310, nx324, nx338, nx352, nx366, nx380, nx394, nx408, nx422, 
      nx432, nx466, nx484, nx496, nx504, nx514, MISR_out_29, MAC0_adderB_28, 
      LFSROUT_17, LFSROUT_18, LFSROUT_19, LFSROUT_20, LFSROUT_21, LFSROUT_22, 
      LFSROUT_23, LFSROUT_24, LFSROUT_25, LFSROUT_26, LFSROUT_27, LFSROUT_28, 
      LFSROUT_29, LFSROUT_30, LFSROUT_31, LFSROUT_0, LFSROUT_1, LFSROUT_2, 
      LFSROUT_3, LFSROUT_4, LFSROUT_5, LFSROUT_6, LFSROUT_7, LFSROUT_8, 
      LFSROUT_9, LFSROUT_10, LFSROUT_11, LFSROUT_12, LFSROUT_13, LFSROUT_14, 
      LFSROUT_15, LFSROUT_16, nx616, nx622, nx644, nx660, nx672, 
      MAC0_MultA_0, nx686, MAC0_MultB_0, nx698, nx704, nx714, nx732, nx740, 
      nx748, nx758, nx768, nx770, nx780, nx788, nx796, nx804, nx814, nx824, 
      nx826, nx828, nx830, nx840, nx848, nx856, nx864, nx872, nx882, nx892, 
      nx894, nx896, nx898, nx900, nx902, nx912, nx920, nx928, nx936, nx944, 
      nx952, nx962, nx972, nx974, nx976, nx978, nx980, nx982, nx984, nx986, 
      nx996, nx1004, nx1012, nx1020, nx1028, nx1036, nx1044, nx1054, nx1064, 
      nx1066, nx1068, nx1070, nx1072, nx1074, nx1076, nx1078, nx1080, nx1082, 
      nx1092, nx1100, nx1108, nx1116, nx1124, nx1132, nx1140, nx1148, nx1158, 
      nx1168, nx1170, nx1172, nx1174, nx1176, nx1178, nx1180, nx1182, nx1184, 
      nx1186, nx1188, nx1190, nx1200, nx1208, nx1216, nx1224, nx1232, nx1240, 
      nx1248, nx1256, nx1264, nx1274, nx1284, nx1286, nx1288, nx1290, nx1292, 
      nx1294, nx1296, nx1298, nx1300, nx1302, nx1304, nx1306, nx1308, nx1310, 
      nx1320, nx1328, nx1336, nx1344, nx1352, nx1360, nx1368, nx1376, nx1384, 
      nx1392, nx1402, nx1412, nx1414, nx1416, nx1418, nx1420, nx1422, nx1424, 
      nx1426, nx1428, nx1430, nx1432, nx1434, nx1436, nx1438, nx1440, nx1442, 
      nx1452, nx1460, nx1468, nx1476, nx1484, nx1492, nx1500, nx1508, nx1516, 
      nx1524, nx1532, nx1542, nx1552, nx1554, nx1556, nx1558, nx1560, nx1562, 
      nx1564, nx1566, nx1568, nx1570, nx1572, nx1574, nx1576, nx1578, nx1580, 
      nx1582, nx1584, nx1586, nx1596, nx1604, nx1612, nx1620, nx1628, nx1636, 
      nx1644, nx1652, nx1660, nx1668, nx1676, nx1684, nx1694, nx1704, nx1706, 
      nx1708, nx1710, nx1712, nx1714, nx1716, nx1718, nx1720, nx1722, nx1724, 
      nx1726, nx1728, nx1730, nx1732, nx1734, nx1736, nx1738, nx1740, nx1742, 
      nx1752, nx1760, nx1768, nx1776, nx1784, nx1792, nx1800, nx1808, nx1816, 
      nx1824, nx1832, nx1840, nx1848, nx1858, nx1868, nx1870, nx1872, nx1874, 
      nx1876, nx1878, nx1880, nx1882, nx1884, nx1886, nx1888, nx1890, nx1892, 
      nx1894, nx1896, nx1898, nx1900, nx1902, nx1904, nx1906, nx1908, nx1910, 
      nx1920, nx1928, nx1936, nx1944, nx1952, nx1960, nx1968, nx1976, nx1984, 
      nx1992, nx2000, nx2008, nx2016, nx2024, nx2034, nx2044, nx2046, nx2048, 
      nx2050, nx2052, nx2054, nx2056, nx2058, nx2060, nx2062, nx2064, nx2066, 
      nx2068, nx2070, nx2072, nx2074, nx2076, nx2078, nx2080, nx2082, nx2084, 
      nx2086, nx2088, nx2090, nx2100, nx2108, nx2116, nx2124, nx2132, nx2140, 
      nx2148, nx2156, nx2164, nx2172, nx2180, nx2188, nx2196, nx2204, nx2212, 
      nx2222, nx2232, nx2234, nx2236, nx2238, nx2240, nx2242, nx2244, nx2246, 
      nx2248, nx2250, nx2252, nx2254, nx2256, nx2258, nx2260, nx2262, nx2264, 
      nx2266, nx2268, nx2270, nx2272, nx2274, nx2276, nx2278, nx2280, nx2282, 
      nx2292, nx2300, nx2412, nx2414, nx2484, nx2492, nx2500, nx2508, nx2516, 
      nx2524, nx2532, nx2540, nx2548, nx2556, nx2564, nx2572, nx2580, nx2588, 
      nx2594, nx2596, nx2602, nx2604, nx2610, nx2612, nx2618, nx2620, nx2626, 
      nx2628, nx2634, nx2636, nx2642, nx2644, nx2650, nx2658, nx2674, nx2682, 
      nx2690, nx2706, nx2714, nx2722, nx2738, nx2746, nx2754, nx2756, nx2758, 
      nx2760, nx2770, nx2772, nx2774, nx2776, nx2786, nx2788, nx2790, nx2792, 
      nx2802, nx2804, nx2818, nx2826, nx2850, nx2858, nx2882, nx2890, nx2914, 
      nx2916, nx2930, nx2932, nx2946, nx2948, nx2958, nx2974, nx2982, nx2990, 
      nx2998, nx3006, nx3014, nx3022, nx3038, nx3046, nx3048, nx3058, nx3060, 
      nx3066, nx3068, nx3070, nx3072, nx3078, nx3080, nx3094, nx3102, nx3118, 
      nx3126, nx3134, nx3142, nx3158, nx3166, nx3178, nx3180, nx3190, nx3192, 
      nx3194, nx3196, nx3198, nx3200, nx3210, nx3212, nx3218, nx3226, nx3234, 
      nx3242, nx3250, nx3258, nx3266, nx3274, nx3282, nx3290, nx3292, nx3294, 
      nx3296, nx3302, nx3304, nx3306, nx3308, nx3310, nx3312, nx3314, nx3316, 
      nx3322, nx3324, nx3338, nx3346, nx3354, nx3362, nx3370, nx3378, nx3402, 
      nx3404, nx3406, nx3408, nx3410, nx3412, nx3414, nx3416, nx3418, nx3420, 
      nx3430, nx3478, nx3486, nx3488, nx3518, nx3526, nx3534, nx3542, nx3550, 
      nx3558, nx3570, nx3572, nx3578, nx3580, nx3586, nx3588, nx3594, nx3602, 
      nx3618, nx3626, nx3634, nx3636, nx3638, nx3640, nx3650, nx3652, nx3666, 
      nx3674, nx3698, nx3700, nx3710, nx3726, nx3734, nx3736, nx3746, 
      MAC0_adderB_27, nx3752, MAC0_adderB_26, nx3758, MAC0_adderB_25, nx3764, 
      MAC0_adderB_24, nx3770, MAC0_adderB_23, nx3776, MAC0_adderB_22, nx3782, 
      MAC0_adderB_21, nx3788, MAC0_adderB_20, nx3794, MAC0_adderB_19, nx3800, 
      MAC0_adderB_18, nx3806, MAC0_adderB_17, nx3812, MAC0_adderB_16, nx3818, 
      MAC0_adderB_15, nx3824, nx3830, MAC0_adderB_14, nx3836, nx3842, 
      MAC0_adderB_13, nx3848, nx3854, MAC0_adderB_12, nx3860, nx3866, 
      MAC0_adderB_11, nx3872, nx3878, MAC0_adderB_10, nx3884, nx3890, 
      MAC0_adderB_9, nx3896, nx3902, MAC0_adderB_8, nx3908, nx3914, 
      MAC0_adderB_7, nx3920, nx3926, MAC0_adderB_6, nx3932, nx3938, 
      MAC0_adderB_5, nx3950, MAC0_adderB_4, nx3962, MAC0_adderB_3, nx3974, 
      MAC0_adderB_2, nx3986, MAC0_adderB_1, nx4000, MAC0_adderB_0, nx989, 
      nx991, nx4040, nx993, nx4046, nx4056, nx995, nx4062, nx4072, nx997, 
      nx4078, nx4088, nx998, nx4094, nx4104, nx999, nx4110, nx4120, nx1000, 
      nx4126, nx4136, nx1001, nx4142, nx4152, nx1003, nx4158, nx4168, nx1005, 
      nx4174, nx4184, nx1007, nx4190, nx4200, nx1009, nx4206, nx4216, nx1011, 
      nx4222, nx4232, nx1013, nx4238, nx4248, nx1015, nx4254, nx4264, nx1017, 
      nx4270, nx4280, nx1019, nx4286, nx4296, nx1021, nx4302, nx4312, nx1023, 
      nx4318, nx4328, nx1025, nx4334, nx4344, nx1027, nx4350, nx4360, nx1029, 
      nx4366, nx4376, nx1031, nx4382, nx4392, nx1033, nx4398, nx4408, nx1035, 
      nx4414, nx4424, nx1037, nx4430, nx4440, nx1039, nx4446, nx4456, nx1041, 
      nx4462, nx4472, MAC0_adderB_29, nx4478, nx4486, nx4498, nx4500, nx4502, 
      nx4508, nx4510, MISR_out_30, nx4522, MAC0_adderB_30, nx4536, nx4538, 
      nx4540, nx4546, nx4548, MISR_out_31, MAC0_adderB_31, nx4566, nx4574, 
      MISR_out_0, MISR_out_1, MISR_out_2, MISR_out_3, MISR_out_4, MISR_out_5, 
      MISR_out_6, MISR_out_7, MISR_out_8, MISR_out_9, MISR_out_10, 
      MISR_out_11, MISR_out_12, MISR_out_13, MISR_out_14, MISR_out_15, 
      MISR_out_16, MISR_out_17, MISR_out_18, MISR_out_19, MISR_out_20, 
      MISR_out_21, MISR_out_22, MISR_out_23, MISR_out_24, MISR_out_25, 
      MISR_out_26, MISR_out_27, MISR_out_28, nx4580, nx4586, nx4592, nx4600, 
      nx4608, nx4614, nx4620, nx4626, nx4632, nx4640, nx4646, nx4652, nx4658, 
      nx4664, nx4670, nx4676, nx4682, nx4688, nx4694, nx4700, nx4706, nx4712, 
      nx4718, nx4724, nx4730, nx4736, nx4742, nx4748, nx4754, nx4760, nx4766, 
      nx4772, nx4784, nx4800, nx4838, nx4848, nx4860, nx4870, nx4876, nx4878, 
      nx1049, nx1059, nx1069, nx1079, nx1089, nx1099, nx1109, nx1119, nx1129, 
      nx1139, nx1149, nx1159, nx1169, nx1179, nx1189, nx1199, nx1209, nx1219, 
      nx1229, nx1239, nx1249, nx1259, nx1269, nx1279, nx1289, nx1299, nx1309, 
      nx1319, nx1329, nx1339, nx1349, nx1359, nx1369, nx1379, nx1389, nx1399, 
      nx1409, nx1419, nx1429, nx1439, nx1449, nx1459, nx1469, nx1479, nx1489, 
      nx1499, nx1509, nx1519, nx1529, nx1539, nx1549, nx1559, nx1569, nx1579, 
      nx1589, nx1599, nx1609, nx1619, nx1629, nx1639, nx1649, nx1659, nx1669, 
      nx1679, nx1689, nx1699, nx1709, nx1719, nx1729, nx1739, nx1749, nx1759, 
      nx1769, nx1779, nx1789, nx1799, nx1809, nx1819, nx1829, nx1839, nx1849, 
      nx1859, nx1869, nx1879, nx1889, nx1899, nx1909, nx1919, nx1929, nx1939, 
      nx1949, nx1959, nx1969, nx1979, nx1989, nx1999, nx2009, nx2019, nx2029, 
      nx2039, nx2049, nx2059, nx2069, nx2079, nx2089, nx2099, nx2109, nx2119, 
      nx2129, nx2139, nx2149, nx2159, nx2169, nx2179, nx2189, nx2199, nx2209, 
      nx2219, nx2229, nx2239, nx2249, nx2259, nx2269, nx2279, nx2289, nx2299, 
      nx2309, nx2319, nx2335, nx2339, nx2347, nx2349, nx2353, nx2359, nx2361, 
      nx2379, nx2389, nx2397, nx2407, nx2413, nx2415, nx2427, nx2433, nx2437, 
      nx2447, nx2453, nx2455, nx2457, nx2467, nx2473, nx2475, nx2485, nx2491, 
      nx2493, nx2497, nx2507, nx2513, nx2515, nx2525, nx2531, nx2533, nx2535, 
      nx2545, nx2551, nx2553, nx2563, nx2569, nx2571, nx2573, nx2583, nx2589, 
      nx2591, nx2601, nx2607, nx2609, nx2611, nx2621, nx2627, nx2629, nx2639, 
      nx2645, nx2655, nx2671, nx2679, nx2687, nx2695, nx2703, nx2711, nx2719, 
      nx2727, nx2735, nx2743, nx2751, nx2759, nx2767, nx2775, nx2783, nx2791, 
      nx2799, nx2807, nx2815, nx2823, nx2831, nx2839, nx2847, nx2855, nx2863, 
      nx2871, nx2879, nx2887, nx2901, nx3115, nx3117, nx3125, nx3131, nx3135, 
      nx3137, nx3143, nx3145, nx3153, nx3159, nx3161, nx3163, nx3165, nx3167, 
      nx3173, nx3179, nx3189, nx3195, nx3197, nx3201, nx3207, nx3209, nx3211, 
      nx3213, nx3219, nx3225, nx3235, nx3241, nx3243, nx3247, nx3251, nx3255, 
      nx3261, nx3263, nx3265, nx3267, nx3273, nx3279, nx3289, nx3295, nx3297, 
      nx3301, nx3305, nx3309, nx3313, nx3319, nx3325, nx3331, nx3333, nx3335, 
      nx3341, nx3347, nx3357, nx3363, nx3365, nx3369, nx3373, nx3377, nx3381, 
      nx3387, nx3391, nx3397, nx3403, nx3409, nx3411, nx3413, nx3419, nx3425, 
      nx3435, nx3441, nx3443, nx3449, nx3453, nx3457, nx3461, nx3467, nx3471, 
      nx3477, nx3481, nx3487, nx3493, nx3499, nx3501, nx3503, nx3509, nx3515, 
      nx3525, nx3531, nx3533, nx3539, nx3543, nx3547, nx3551, nx3557, nx3561, 
      nx3567, nx3571, nx3577, nx3581, nx3587, nx3593, nx3599, nx3601, nx3603, 
      nx3609, nx3615, nx3625, nx3631, nx3633, nx3639, nx3643, nx3647, nx3651, 
      nx3657, nx3661, nx3667, nx3671, nx3677, nx3681, nx3687, nx3691, nx3697, 
      nx3703, nx3709, nx3711, nx3713, nx3719, nx3725, nx3735, nx3741, nx3743, 
      nx3749, nx3753, nx3756, nx3759, nx3763, nx3767, nx3771, nx3774, nx3779, 
      nx3783, nx3787, nx3791, nx3795, nx3798, nx3803, nx3807, nx3811, nx3813, 
      nx3815, nx3819, nx3823, nx3833, nx3837, nx3839, nx3845, nx3849, nx3853, 
      nx3857, nx3861, nx3865, nx3870, nx3873, nx3879, nx3882, nx3887, nx3891, 
      nx3895, nx3899, nx3905, nx3909, nx3915, nx3919, nx3925, nx3927, nx3929, 
      nx3933, nx3939, nx3947, nx3953, nx3955, nx3961, nx3965, nx3969, nx3973, 
      nx3978, nx3981, nx3987, nx3990, nx3995, nx3999, nx4004, nx4007, nx4011, 
      nx4015, nx4019, nx4023, nx4027, nx4031, nx4037, nx4043, nx4047, nx4049, 
      nx4051, nx4057, nx4061, nx4071, nx4076, nx4079, nx4085, nx4089, nx4092, 
      nx4095, nx4101, nx4105, nx4109, nx4113, nx4119, nx4123, nx4127, nx4131, 
      nx4137, nx4140, nx4145, nx4149, nx4155, nx4159, nx4165, nx4169, nx4173, 
      nx4179, nx4185, nx4187, nx4189, nx4195, nx4201, nx4209, nx4215, nx4217, 
      nx4221, nx4225, nx4229, nx4233, nx4237, nx4241, nx4247, nx4251, nx4255, 
      nx4259, nx4265, nx4268, nx4273, nx4277, nx4283, nx4287, nx4293, nx4297, 
      nx4301, nx4305, nx4311, nx4315, nx4319, nx4325, nx4331, nx4333, nx4335, 
      nx4341, nx4347, nx4357, nx4363, nx4365, nx4371, nx4375, nx4379, nx4383, 
      nx4389, nx4393, nx4397, nx4401, nx4407, nx4411, nx4415, nx4419, nx4425, 
      nx4428, nx4433, nx4437, nx4443, nx4447, nx4453, nx4457, nx4461, nx4465, 
      nx4471, nx4475, nx4481, nx4487, nx4493, nx4495, nx4497, nx4503, nx4507, 
      nx4516, nx4519, nx4521, nx4523, nx4525, nx4527, nx4529, nx4531, nx4535, 
      nx4537, nx4539, nx4541, nx4544, nx4547, nx4549, nx4551, nx4554, nx4557, 
      nx4559, nx4561, nx4565, nx4567, nx4569, nx4571, nx4575, nx4577, nx4579, 
      nx4581, nx4584, nx4587, nx4589, nx4591, nx4595, nx4597, nx4599, nx4601, 
      nx4604, nx4607, nx4609, nx4611, nx4615, nx4617, nx4619, nx4621, nx4624, 
      nx4627, nx4629, nx4631, nx4635, nx4637, nx4639, nx4641, nx4644, nx4647, 
      nx4649, nx4651, nx4656, nx4665, nx4674, nx4677, nx4681, nx4683, nx4685, 
      nx4689, nx4693, nx4695, nx4697, nx4701, nx4705, nx4707, nx4709, nx4713, 
      nx4717, nx4719, nx4721, nx4725, nx4729, nx4731, nx4733, nx4737, nx4741, 
      nx4743, nx4745, nx4749, nx4753, nx4755, nx4757, nx4763, nx4771, nx4775, 
      nx4779, nx4781, nx4783, nx4785, nx4787, nx4789, nx4791, nx4793, nx4797, 
      nx4801, nx4805, nx4809, nx4815, nx4817, nx4819, nx4821, nx4823, nx4825, 
      nx4827, nx4829, nx4833, nx4837, nx4841, nx4845, nx4851, nx4853, nx4855, 
      nx4857, nx4859, nx4861, nx4863, nx4865, nx4869, nx4873, nx4877, nx4881, 
      nx4884, nx4889, nx4896, nx4899, nx4901, nx4903, nx4906, nx4911, nx4915, 
      nx4917, nx4919, nx4921, nx4923, nx4925, nx4927, nx4929, nx4932, nx4934, 
      nx4936, nx4939, nx4944, nx4948, nx4950, nx4952, nx4954, nx4956, nx4958, 
      nx4960, nx4962, nx4965, nx4967, nx4969, nx4972, nx4977, nx4981, nx4983, 
      nx4985, nx4987, nx4989, nx4991, nx4993, nx4999, nx5007, nx5009, nx5011, 
      nx5013, nx5015, nx5017, nx5019, nx5022, nx5025, nx5029, nx5031, nx5033, 
      nx5037, nx5040, nx5043, nx5047, nx5049, nx5051, nx5053, nx5057, nx5061, 
      nx5063, nx5065, nx5067, nx5069, nx5071, nx5073, nx5076, nx5079, nx5085, 
      nx5093, nx5096, nx5100, nx5102, nx5104, nx5106, nx5108, nx5110, nx5112, 
      nx5115, nx5118, nx5121, nx5124, nx5127, nx5131, nx5135, nx5139, nx5141, 
      nx5143, nx5145, nx5147, nx5149, nx5151, nx5154, nx5157, nx5161, nx5163, 
      nx5165, nx5170, nx5177, nx5180, nx5184, nx5186, nx5188, nx5190, nx5194, 
      nx5197, nx5200, nx5203, nx5207, nx5210, nx5214, nx5218, nx5222, nx5224, 
      nx5226, nx5230, nx5233, nx5236, nx5239, nx5244, nx5251, nx5254, nx5256, 
      nx5258, nx5261, nx5266, nx5269, nx5272, nx5275, nx5279, nx5282, nx5286, 
      nx5289, nx5293, nx5297, nx5301, nx5303, nx5305, nx5307, nx5309, nx5311, 
      nx5313, nx5319, nx5327, nx5329, nx5331, nx5333, nx5335, nx5337, nx5339, 
      nx5341, nx5344, nx5346, nx5348, nx5350, nx5353, nx5355, nx5357, nx5359, 
      nx5362, nx5364, nx5366, nx5368, nx5371, nx5373, nx5375, nx5378, nx5383, 
      nx5389, nx5397, nx5400, nx5404, nx5406, nx5408, nx5412, nx5416, nx5418, 
      nx5420, nx5424, nx5428, nx5430, nx5432, nx5437, nx5444, nx5447, nx5451, 
      nx5453, nx5455, nx5457, nx5459, nx5461, nx5463, nx5465, nx5468, nx5471, 
      nx5474, nx5477, nx5480, nx5485, nx5492, nx5495, nx5497, nx5499, nx5502, 
      nx5507, nx5511, nx5513, nx5515, nx5517, nx5519, nx5521, nx5523, nx5529, 
      nx5537, nx5539, nx5541, nx5543, nx5545, nx5547, nx5549, nx5552, nx5555, 
      nx5561, nx5569, nx5572, nx5576, nx5578, nx5580, nx5584, nx5592, nx5595, 
      nx5602, nx5605, nx5608, nx5620, nx5623, nx5626, nx5633, nx5638, nx5643, 
      nx5648, nx5653, nx5678, nx5683, nx5688, nx5693, nx5698, nx5703, nx5708, 
      nx5713, nx5718, nx5723, nx5728, nx5733, nx5738, nx5743, nx5753, nx5758, 
      nx5763, nx5773, nx5778, nx5780, nx5782, nx5784, nx5786, nx5788, nx5800, 
      nx5802, nx5804, nx5806, nx5808, nx5810, nx5812, nx5814, nx5816, nx5818, 
      nx5820, nx5822, nx5824, nx5844, nx5848, nx5850, nx5852, nx5854, nx5856, 
      nx5860, nx5862, nx5864, nx5866, nx5868, nx5870, nx5872, nx5874, nx5876, 
      nx5878, nx5880, nx5882, nx5884, nx5886, nx5888, nx5890, nx5892, nx5894, 
      nx5896, nx5898, nx5900, nx5902, nx5904, nx5906, nx5908, nx5910, nx5912, 
      nx5914, nx5916, nx5918, nx5920, nx5922, nx5924, nx5926, nx5928, nx5930, 
      nx5932, nx5934, nx5936, nx5938, nx5940, nx5942, nx5944, nx5946, nx5948, 
      nx5950, nx5952, nx5954, nx5956, nx5958, nx5960, nx5962, nx5964, nx5966, 
      nx5968, nx5970, nx5972, nx5974, nx5980, nx5982, nx5984, nx5986, nx5988, 
      nx5990, nx5992, nx5994, nx5996, nx5998, nx6000, nx6002, nx6004, nx6006, 
      nx6008, nx6010, nx6012, nx6014, nx6016, nx6018, nx6020, nx6022, nx6024, 
      nx6026, nx6028, nx6030, nx6032, nx6034, nx6036, nx6038, nx6040, nx6042, 
      nx6044, nx6046, nx6048, nx6050, nx6052, nx6054, nx6056, nx6058, nx6060, 
      nx6062, nx6064, nx6066, nx6068, nx6070, nx6072, nx6074, nx6076, nx6078, 
      nx6080, nx6082, nx6084, nx6086, nx6088, nx6090, nx6092, nx6094, nx6096, 
      nx6098, nx6100, nx6102, nx6104, nx6106, nx6108, nx6110, nx6112, nx6114, 
      nx6116, nx6118, nx6120, nx6122, nx6124, nx6126, nx6128, nx6130, nx6132, 
      nx6134, nx6136, nx6138, nx6140: std_logic ;

begin
   RegOut(31) <= RegOut_dup0_31 ;
   RegOut(30) <= RegOut_dup0_30 ;
   RegOut(29) <= RegOut_dup0_29 ;
   RegOut(28) <= RegOut_dup0_28 ;
   RegOut(27) <= RegOut_dup0_27 ;
   RegOut(26) <= RegOut_dup0_26 ;
   RegOut(25) <= RegOut_dup0_25 ;
   RegOut(24) <= RegOut_dup0_24 ;
   RegOut(23) <= RegOut_dup0_23 ;
   RegOut(22) <= RegOut_dup0_22 ;
   RegOut(21) <= RegOut_dup0_21 ;
   RegOut(20) <= RegOut_dup0_20 ;
   RegOut(19) <= RegOut_dup0_19 ;
   RegOut(18) <= RegOut_dup0_18 ;
   RegOut(17) <= RegOut_dup0_17 ;
   RegOut(16) <= RegOut_dup0_16 ;
   RegOut(15) <= RegOut_dup0_15 ;
   RegOut(14) <= RegOut_dup0_14 ;
   RegOut(13) <= RegOut_dup0_13 ;
   RegOut(12) <= RegOut_dup0_12 ;
   RegOut(11) <= RegOut_dup0_11 ;
   RegOut(10) <= RegOut_dup0_10 ;
   RegOut(9) <= RegOut_dup0_9 ;
   RegOut(8) <= RegOut_dup0_8 ;
   RegOut(7) <= RegOut_dup0_7 ;
   RegOut(6) <= RegOut_dup0_6 ;
   RegOut(5) <= RegOut_dup0_5 ;
   RegOut(4) <= RegOut_dup0_4 ;
   RegOut(3) <= RegOut_dup0_3 ;
   RegOut(2) <= RegOut_dup0_2 ;
   RegOut(1) <= RegOut_dup0_1 ;
   RegOut(0) <= RegOut_dup0_0 ;
   Pass <= Pass_dup0 ;
   Complete <= Complete_dup0 ;
   TEST0_reg_complete_v : dffr port map ( Q=>Complete_dup0, QB=>OPEN, D=>
      nx514, CLK=>clk, R=>nx5804);
   ix515 : or02 port map ( Y=>nx514, A0=>nx2335, A1=>Complete_dup0);
   ix2336 : nor04 port map ( Y=>nx2335, A0=>nx504, A1=>nx496, A2=>nx484, A3
      =>nx466);
   COUNT0_REG0_reg_Y_0 : dffr port map ( Q=>CounterOut_0, QB=>nx2339, D=>
      nx1049, CLK=>clk, R=>nx5800);
   TEST0_reg_TestEN : dffr port map ( Q=>OPEN, QB=>nx2347, D=>StartTest, CLK
      =>clk, R=>nx5800);
   ix1060 : oai21 port map ( Y=>nx1059, A0=>nx2353, A1=>nx5998, B0=>nx2359);
   ix2354 : oai21 port map ( Y=>nx2353, A0=>CounterOut_0, A1=>CounterOut_1, 
      B0=>nx987);
   COUNT0_REG0_reg_Y_1 : dffr port map ( Q=>CounterOut_1, QB=>nx2349, D=>
      nx1059, CLK=>clk, R=>nx5800);
   ix2360 : nand02 port map ( Y=>nx2359, A0=>CounterOut_1, A1=>nx5998);
   COUNT0_REG0_reg_Y_2 : dffr port map ( Q=>CounterOut_2, QB=>nx2361, D=>
      nx1069, CLK=>clk, R=>nx5800);
   COUNT0_REG0_reg_Y_3 : dffr port map ( Q=>CounterOut_3, QB=>OPEN, D=>
      nx1079, CLK=>clk, R=>nx5800);
   ix45 : xnor2 port map ( Y=>nx44, A0=>nx985, A1=>CounterOut_3);
   COUNT0_REG0_reg_Y_4 : dffr port map ( Q=>CounterOut_4, QB=>nx2379, D=>
      nx1089, CLK=>clk, R=>nx5800);
   ix59 : aoi21 port map ( Y=>nx58, A0=>nx983, A1=>nx2379, B0=>nx2389);
   COUNT0_REG0_reg_Y_5 : dffr port map ( Q=>CounterOut_5, QB=>nx2397, D=>
      nx1099, CLK=>clk, R=>nx5800);
   COUNT0_REG0_reg_Y_6 : dffr port map ( Q=>CounterOut_6, QB=>nx2407, D=>
      nx1109, CLK=>clk, R=>nx5800);
   ix81 : nand02 port map ( Y=>nx979, A0=>nx2389, A1=>CounterOut_5);
   COUNT0_REG0_reg_Y_7 : dffr port map ( Q=>CounterOut_7, QB=>nx2415, D=>
      nx1119, CLK=>clk, R=>nx5800);
   ix485 : nand04 port map ( Y=>nx484, A0=>CounterOut_8, A1=>CounterOut_9, 
      A2=>nx2437, A3=>nx2457);
   COUNT0_REG0_reg_Y_8 : dffr port map ( Q=>CounterOut_8, QB=>nx2427, D=>
      nx1129, CLK=>clk, R=>nx5800);
   ix109 : nand02 port map ( Y=>nx975, A0=>nx2413, A1=>CounterOut_7);
   COUNT0_REG0_reg_Y_9 : dffr port map ( Q=>CounterOut_9, QB=>OPEN, D=>
      nx1139, CLK=>clk, R=>nx5800);
   COUNT0_REG0_reg_Y_10 : dffr port map ( Q=>CounterOut_10, QB=>nx2447, D=>
      nx1149, CLK=>clk, R=>nx5800);
   ix137 : nand02 port map ( Y=>nx971, A0=>nx2433, A1=>CounterOut_9);
   COUNT0_REG0_reg_Y_11 : dffr port map ( Q=>CounterOut_11, QB=>nx2455, D=>
      nx1159, CLK=>clk, R=>nx5800);
   COUNT0_REG0_reg_Y_12 : dffr port map ( Q=>CounterOut_12, QB=>nx2467, D=>
      nx1169, CLK=>clk, R=>nx5800);
   ix165 : nand02 port map ( Y=>nx967, A0=>nx2453, A1=>CounterOut_11);
   COUNT0_REG0_reg_Y_13 : dffr port map ( Q=>CounterOut_13, QB=>nx2475, D=>
      nx1179, CLK=>clk, R=>nx5800);
   COUNT0_REG0_reg_Y_14 : dffr port map ( Q=>CounterOut_14, QB=>nx2485, D=>
      nx1189, CLK=>clk, R=>nx5802);
   ix193 : nand02 port map ( Y=>nx965, A0=>nx2473, A1=>CounterOut_13);
   COUNT0_REG0_reg_Y_15 : dffr port map ( Q=>CounterOut_15, QB=>nx2493, D=>
      nx1199, CLK=>clk, R=>nx5802);
   ix467 : nand04 port map ( Y=>nx466, A0=>nx2497, A1=>nx2535, A2=>nx2573, 
      A3=>nx2611);
   COUNT0_REG0_reg_Y_16 : dffr port map ( Q=>CounterOut_16, QB=>nx2507, D=>
      nx1209, CLK=>clk, R=>nx5802);
   ix221 : nand02 port map ( Y=>nx963, A0=>nx2491, A1=>CounterOut_15);
   COUNT0_REG0_reg_Y_17 : dffr port map ( Q=>CounterOut_17, QB=>nx2515, D=>
      nx1219, CLK=>clk, R=>nx5802);
   COUNT0_REG0_reg_Y_18 : dffr port map ( Q=>CounterOut_18, QB=>nx2525, D=>
      nx1229, CLK=>clk, R=>nx5802);
   ix249 : nand02 port map ( Y=>nx959, A0=>nx2513, A1=>CounterOut_17);
   COUNT0_REG0_reg_Y_19 : dffr port map ( Q=>CounterOut_19, QB=>nx2533, D=>
      nx1239, CLK=>clk, R=>nx5802);
   COUNT0_REG0_reg_Y_20 : dffr port map ( Q=>CounterOut_20, QB=>nx2545, D=>
      nx1249, CLK=>clk, R=>nx5802);
   ix277 : nand02 port map ( Y=>nx955, A0=>nx2531, A1=>CounterOut_19);
   COUNT0_REG0_reg_Y_21 : dffr port map ( Q=>CounterOut_21, QB=>nx2553, D=>
      nx1259, CLK=>clk, R=>nx5802);
   COUNT0_REG0_reg_Y_22 : dffr port map ( Q=>CounterOut_22, QB=>nx2563, D=>
      nx1269, CLK=>clk, R=>nx5802);
   ix305 : nand02 port map ( Y=>nx951, A0=>nx2551, A1=>CounterOut_21);
   COUNT0_REG0_reg_Y_23 : dffr port map ( Q=>CounterOut_23, QB=>nx2571, D=>
      nx1279, CLK=>clk, R=>nx5802);
   COUNT0_REG0_reg_Y_24 : dffr port map ( Q=>CounterOut_24, QB=>nx2583, D=>
      nx1289, CLK=>clk, R=>nx5802);
   ix333 : nand02 port map ( Y=>nx947, A0=>nx2569, A1=>CounterOut_23);
   COUNT0_REG0_reg_Y_25 : dffr port map ( Q=>CounterOut_25, QB=>nx2591, D=>
      nx1299, CLK=>clk, R=>nx5802);
   COUNT0_REG0_reg_Y_26 : dffr port map ( Q=>CounterOut_26, QB=>nx2601, D=>
      nx1309, CLK=>clk, R=>nx5802);
   ix361 : nand02 port map ( Y=>nx943, A0=>nx2589, A1=>CounterOut_25);
   COUNT0_REG0_reg_Y_27 : dffr port map ( Q=>CounterOut_27, QB=>nx2609, D=>
      nx1319, CLK=>clk, R=>nx5802);
   COUNT0_REG0_reg_Y_28 : dffr port map ( Q=>CounterOut_28, QB=>nx2621, D=>
      nx1329, CLK=>clk, R=>nx5802);
   ix389 : nand02 port map ( Y=>nx939, A0=>nx2607, A1=>CounterOut_27);
   COUNT0_REG0_reg_Y_29 : dffr port map ( Q=>CounterOut_29, QB=>nx2629, D=>
      nx1339, CLK=>clk, R=>nx5804);
   COUNT0_REG0_reg_Y_30 : dffr port map ( Q=>CounterOut_30, QB=>nx2639, D=>
      nx1349, CLK=>clk, R=>nx5804);
   ix417 : nand02 port map ( Y=>nx935, A0=>nx2627, A1=>CounterOut_29);
   COUNT0_REG0_reg_Y_31 : dffr port map ( Q=>CounterOut_31, QB=>OPEN, D=>
      nx1359, CLK=>clk, R=>nx5804);
   ix433 : xor2 port map ( Y=>nx432, A0=>CounterOut_31, A1=>nx2645);
   TEST0_reg_pass_v : dffr port map ( Q=>Pass_dup0, QB=>OPEN, D=>nx4878, CLK
      =>clk, R=>nx5824);
   ix4879 : or02 port map ( Y=>nx4878, A0=>nx4876, A1=>Pass_dup0);
   ix4877 : nor04 port map ( Y=>nx4876, A0=>nx2655, A1=>nx5784, A2=>nx5786, 
      A3=>nx5788);
   ix2656 : nand04 port map ( Y=>nx2655, A0=>nx4784, A1=>nx5773, A2=>
      MISR_out_27, A3=>nx4800);
   MAC0_BigBoyReg_reg_Y_29 : dffr port map ( Q=>RegOut_dup0_29, QB=>OPEN, D
      =>nx1979, CLK=>clk, R=>nx5820);
   ix1980 : mux21 port map ( Y=>nx1979, A0=>RegOut_dup0_29, A1=>nx4510, S0=>
      WE);
   ix2672 : aoi22 port map ( Y=>nx2671, A0=>RegOut_dup0_28, A1=>nx4456, B0=>
      MAC0_adderB_28, B1=>nx5561);
   MAC0_BigBoyReg_reg_Y_28 : dffr port map ( Q=>RegOut_dup0_28, QB=>OPEN, D
      =>nx1969, CLK=>clk, R=>nx5820);
   ix1970 : mux21 port map ( Y=>nx1969, A0=>RegOut_dup0_28, A1=>nx1041, S0=>
      WE);
   ix2680 : aoi22 port map ( Y=>nx2679, A0=>RegOut_dup0_27, A1=>nx4440, B0=>
      MAC0_adderB_27, B1=>nx5529);
   MAC0_BigBoyReg_reg_Y_27 : dffr port map ( Q=>RegOut_dup0_27, QB=>OPEN, D
      =>nx1959, CLK=>clk, R=>nx5820);
   ix1960 : mux21 port map ( Y=>nx1959, A0=>RegOut_dup0_27, A1=>nx1039, S0=>
      WE);
   ix2688 : aoi22 port map ( Y=>nx2687, A0=>RegOut_dup0_26, A1=>nx4424, B0=>
      MAC0_adderB_26, B1=>nx5485);
   MAC0_BigBoyReg_reg_Y_26 : dffr port map ( Q=>RegOut_dup0_26, QB=>OPEN, D
      =>nx1949, CLK=>clk, R=>nx5820);
   ix1950 : mux21 port map ( Y=>nx1949, A0=>RegOut_dup0_26, A1=>nx1037, S0=>
      WE);
   ix2696 : aoi22 port map ( Y=>nx2695, A0=>RegOut_dup0_25, A1=>nx4408, B0=>
      MAC0_adderB_25, B1=>nx5437);
   MAC0_BigBoyReg_reg_Y_25 : dffr port map ( Q=>RegOut_dup0_25, QB=>OPEN, D
      =>nx1939, CLK=>clk, R=>nx5818);
   ix1940 : mux21 port map ( Y=>nx1939, A0=>RegOut_dup0_25, A1=>nx1035, S0=>
      WE);
   ix2704 : aoi22 port map ( Y=>nx2703, A0=>RegOut_dup0_24, A1=>nx4392, B0=>
      MAC0_adderB_24, B1=>nx5389);
   MAC0_BigBoyReg_reg_Y_24 : dffr port map ( Q=>RegOut_dup0_24, QB=>OPEN, D
      =>nx1929, CLK=>clk, R=>nx5818);
   ix1930 : mux21 port map ( Y=>nx1929, A0=>RegOut_dup0_24, A1=>nx1033, S0=>
      WE);
   ix2712 : aoi22 port map ( Y=>nx2711, A0=>RegOut_dup0_23, A1=>nx4376, B0=>
      MAC0_adderB_23, B1=>nx5319);
   MAC0_BigBoyReg_reg_Y_23 : dffr port map ( Q=>RegOut_dup0_23, QB=>OPEN, D
      =>nx1919, CLK=>clk, R=>nx5818);
   ix1920 : mux21 port map ( Y=>nx1919, A0=>RegOut_dup0_23, A1=>nx1031, S0=>
      WE);
   ix2720 : aoi22 port map ( Y=>nx2719, A0=>RegOut_dup0_22, A1=>nx4360, B0=>
      MAC0_adderB_22, B1=>nx5244);
   MAC0_BigBoyReg_reg_Y_22 : dffr port map ( Q=>RegOut_dup0_22, QB=>OPEN, D
      =>nx1909, CLK=>clk, R=>nx5818);
   ix1910 : mux21 port map ( Y=>nx1909, A0=>RegOut_dup0_22, A1=>nx1029, S0=>
      WE);
   ix2728 : aoi22 port map ( Y=>nx2727, A0=>RegOut_dup0_21, A1=>nx4344, B0=>
      MAC0_adderB_21, B1=>nx5170);
   MAC0_BigBoyReg_reg_Y_21 : dffr port map ( Q=>RegOut_dup0_21, QB=>OPEN, D
      =>nx1899, CLK=>clk, R=>nx5818);
   ix1900 : mux21 port map ( Y=>nx1899, A0=>RegOut_dup0_21, A1=>nx1027, S0=>
      WE);
   ix2736 : aoi22 port map ( Y=>nx2735, A0=>RegOut_dup0_20, A1=>nx4328, B0=>
      MAC0_adderB_20, B1=>nx5085);
   MAC0_BigBoyReg_reg_Y_20 : dffr port map ( Q=>RegOut_dup0_20, QB=>OPEN, D
      =>nx1889, CLK=>clk, R=>nx5818);
   ix1890 : mux21 port map ( Y=>nx1889, A0=>RegOut_dup0_20, A1=>nx1025, S0=>
      WE);
   ix2744 : aoi22 port map ( Y=>nx2743, A0=>RegOut_dup0_19, A1=>nx4312, B0=>
      MAC0_adderB_19, B1=>nx4999);
   MAC0_BigBoyReg_reg_Y_19 : dffr port map ( Q=>RegOut_dup0_19, QB=>OPEN, D
      =>nx1879, CLK=>clk, R=>nx5818);
   ix1880 : mux21 port map ( Y=>nx1879, A0=>RegOut_dup0_19, A1=>nx1023, S0=>
      WE);
   ix2752 : aoi22 port map ( Y=>nx2751, A0=>RegOut_dup0_18, A1=>nx4296, B0=>
      MAC0_adderB_18, B1=>nx4889);
   MAC0_BigBoyReg_reg_Y_18 : dffr port map ( Q=>RegOut_dup0_18, QB=>OPEN, D
      =>nx1869, CLK=>clk, R=>nx5818);
   ix1870 : mux21 port map ( Y=>nx1869, A0=>RegOut_dup0_18, A1=>nx1021, S0=>
      WE);
   ix2760 : aoi22 port map ( Y=>nx2759, A0=>RegOut_dup0_17, A1=>nx4280, B0=>
      MAC0_adderB_17, B1=>nx4763);
   MAC0_BigBoyReg_reg_Y_17 : dffr port map ( Q=>RegOut_dup0_17, QB=>OPEN, D
      =>nx1859, CLK=>clk, R=>nx5816);
   ix1860 : mux21 port map ( Y=>nx1859, A0=>RegOut_dup0_17, A1=>nx1019, S0=>
      WE);
   ix2768 : aoi22 port map ( Y=>nx2767, A0=>RegOut_dup0_16, A1=>nx4264, B0=>
      MAC0_adderB_16, B1=>nx4665);
   MAC0_BigBoyReg_reg_Y_16 : dffr port map ( Q=>RegOut_dup0_16, QB=>OPEN, D
      =>nx1849, CLK=>clk, R=>nx5816);
   ix1850 : mux21 port map ( Y=>nx1849, A0=>RegOut_dup0_16, A1=>nx1017, S0=>
      WE);
   ix2776 : aoi22 port map ( Y=>nx2775, A0=>RegOut_dup0_15, A1=>nx4248, B0=>
      MAC0_adderB_15, B1=>nx4507);
   MAC0_BigBoyReg_reg_Y_15 : dffr port map ( Q=>RegOut_dup0_15, QB=>OPEN, D
      =>nx1839, CLK=>clk, R=>nx5816);
   ix1840 : mux21 port map ( Y=>nx1839, A0=>RegOut_dup0_15, A1=>nx1015, S0=>
      WE);
   ix2784 : aoi22 port map ( Y=>nx2783, A0=>RegOut_dup0_14, A1=>nx4232, B0=>
      MAC0_adderB_14, B1=>nx4347);
   MAC0_BigBoyReg_reg_Y_14 : dffr port map ( Q=>RegOut_dup0_14, QB=>OPEN, D
      =>nx1829, CLK=>clk, R=>nx5816);
   ix1830 : mux21 port map ( Y=>nx1829, A0=>RegOut_dup0_14, A1=>nx1013, S0=>
      WE);
   ix2792 : aoi22 port map ( Y=>nx2791, A0=>RegOut_dup0_13, A1=>nx4216, B0=>
      MAC0_adderB_13, B1=>nx4201);
   MAC0_BigBoyReg_reg_Y_13 : dffr port map ( Q=>RegOut_dup0_13, QB=>OPEN, D
      =>nx1819, CLK=>clk, R=>nx5816);
   ix1820 : mux21 port map ( Y=>nx1819, A0=>RegOut_dup0_13, A1=>nx1011, S0=>
      WE);
   ix2800 : aoi22 port map ( Y=>nx2799, A0=>RegOut_dup0_12, A1=>nx4200, B0=>
      MAC0_adderB_12, B1=>nx4061);
   MAC0_BigBoyReg_reg_Y_12 : dffr port map ( Q=>RegOut_dup0_12, QB=>OPEN, D
      =>nx1809, CLK=>clk, R=>nx5814);
   ix1810 : mux21 port map ( Y=>nx1809, A0=>RegOut_dup0_12, A1=>nx1009, S0=>
      WE);
   ix2808 : aoi22 port map ( Y=>nx2807, A0=>RegOut_dup0_11, A1=>nx4184, B0=>
      MAC0_adderB_11, B1=>nx3939);
   MAC0_BigBoyReg_reg_Y_11 : dffr port map ( Q=>RegOut_dup0_11, QB=>OPEN, D
      =>nx1799, CLK=>clk, R=>nx5814);
   ix1800 : mux21 port map ( Y=>nx1799, A0=>RegOut_dup0_11, A1=>nx1007, S0=>
      WE);
   ix2816 : aoi22 port map ( Y=>nx2815, A0=>RegOut_dup0_10, A1=>nx4168, B0=>
      MAC0_adderB_10, B1=>nx3823);
   MAC0_BigBoyReg_reg_Y_10 : dffr port map ( Q=>RegOut_dup0_10, QB=>OPEN, D
      =>nx1789, CLK=>clk, R=>nx5814);
   ix1790 : mux21 port map ( Y=>nx1789, A0=>RegOut_dup0_10, A1=>nx1005, S0=>
      WE);
   ix2824 : aoi22 port map ( Y=>nx2823, A0=>RegOut_dup0_9, A1=>nx4152, B0=>
      MAC0_adderB_9, B1=>nx3725);
   MAC0_BigBoyReg_reg_Y_9 : dffr port map ( Q=>RegOut_dup0_9, QB=>OPEN, D=>
      nx1779, CLK=>clk, R=>nx5814);
   ix1780 : mux21 port map ( Y=>nx1779, A0=>RegOut_dup0_9, A1=>nx1003, S0=>
      WE);
   ix2832 : aoi22 port map ( Y=>nx2831, A0=>RegOut_dup0_8, A1=>nx4136, B0=>
      MAC0_adderB_8, B1=>nx3615);
   MAC0_BigBoyReg_reg_Y_8 : dffr port map ( Q=>RegOut_dup0_8, QB=>OPEN, D=>
      nx1769, CLK=>clk, R=>nx5812);
   ix1770 : mux21 port map ( Y=>nx1769, A0=>RegOut_dup0_8, A1=>nx1001, S0=>
      WE);
   ix2840 : aoi22 port map ( Y=>nx2839, A0=>RegOut_dup0_7, A1=>nx4120, B0=>
      MAC0_adderB_7, B1=>nx3515);
   MAC0_BigBoyReg_reg_Y_7 : dffr port map ( Q=>RegOut_dup0_7, QB=>OPEN, D=>
      nx1759, CLK=>clk, R=>nx5812);
   ix1760 : mux21 port map ( Y=>nx1759, A0=>RegOut_dup0_7, A1=>nx1000, S0=>
      WE);
   ix2848 : aoi22 port map ( Y=>nx2847, A0=>RegOut_dup0_6, A1=>nx4104, B0=>
      MAC0_adderB_6, B1=>nx3425);
   MAC0_BigBoyReg_reg_Y_6 : dffr port map ( Q=>RegOut_dup0_6, QB=>OPEN, D=>
      nx1749, CLK=>clk, R=>nx5812);
   ix1750 : mux21 port map ( Y=>nx1749, A0=>RegOut_dup0_6, A1=>nx999, S0=>WE
   );
   ix2856 : aoi22 port map ( Y=>nx2855, A0=>RegOut_dup0_5, A1=>nx4088, B0=>
      MAC0_adderB_5, B1=>nx3347);
   MAC0_BigBoyReg_reg_Y_5 : dffr port map ( Q=>RegOut_dup0_5, QB=>OPEN, D=>
      nx1739, CLK=>clk, R=>nx5810);
   ix1740 : mux21 port map ( Y=>nx1739, A0=>RegOut_dup0_5, A1=>nx998, S0=>WE
   );
   ix2864 : aoi22 port map ( Y=>nx2863, A0=>RegOut_dup0_4, A1=>nx4072, B0=>
      MAC0_adderB_4, B1=>nx3279);
   MAC0_BigBoyReg_reg_Y_4 : dffr port map ( Q=>RegOut_dup0_4, QB=>OPEN, D=>
      nx1729, CLK=>clk, R=>nx5810);
   ix1730 : mux21 port map ( Y=>nx1729, A0=>RegOut_dup0_4, A1=>nx997, S0=>WE
   );
   ix2872 : aoi22 port map ( Y=>nx2871, A0=>RegOut_dup0_3, A1=>nx4056, B0=>
      MAC0_adderB_3, B1=>nx3225);
   MAC0_BigBoyReg_reg_Y_3 : dffr port map ( Q=>RegOut_dup0_3, QB=>OPEN, D=>
      nx1719, CLK=>clk, R=>nx5810);
   ix1720 : mux21 port map ( Y=>nx1719, A0=>RegOut_dup0_3, A1=>nx995, S0=>WE
   );
   ix2880 : aoi22 port map ( Y=>nx2879, A0=>RegOut_dup0_2, A1=>nx4040, B0=>
      MAC0_adderB_2, B1=>nx3179);
   MAC0_BigBoyReg_reg_Y_2 : dffr port map ( Q=>RegOut_dup0_2, QB=>OPEN, D=>
      nx1709, CLK=>clk, R=>nx5810);
   ix1710 : mux21 port map ( Y=>nx1709, A0=>RegOut_dup0_2, A1=>nx993, S0=>WE
   );
   ix2888 : aoi32 port map ( Y=>nx2887, A0=>RegOut_dup0_1, A1=>RegOut_dup0_0, 
      A2=>MAC0_adderB_0, B0=>MAC0_adderB_1, B1=>nx3143);
   MAC0_BigBoyReg_reg_Y_1 : dffr port map ( Q=>RegOut_dup0_1, QB=>OPEN, D=>
      nx1699, CLK=>clk, R=>nx5808);
   ix1700 : mux21 port map ( Y=>nx1699, A0=>RegOut_dup0_1, A1=>nx991, S0=>WE
   );
   ix4023 : nand02 port map ( Y=>nx989, A0=>RegOut_dup0_0, A1=>MAC0_adderB_0
   );
   MAC0_BigBoyReg_reg_Y_0 : dffr port map ( Q=>RegOut_dup0_0, QB=>OPEN, D=>
      nx1689, CLK=>clk, R=>nx5808);
   ix1690 : oai21 port map ( Y=>nx1689, A0=>nx2901, A1=>nx3115, B0=>nx3117);
   ix2902 : oai21 port map ( Y=>nx2901, A0=>RegOut_dup0_0, A1=>MAC0_adderB_0, 
      B0=>nx989);
   MAC0_RegMultOut_reg_Y_0 : dffr port map ( Q=>MAC0_adderB_0, QB=>OPEN, D=>
      nx704, CLK=>clk, R=>nx5808);
   MAC0_RegMultInA_reg_Y_0 : dffr port map ( Q=>MAC0_MultA_0, QB=>OPEN, D=>
      nx686, CLK=>clk, R=>nx5808);
   LFSR0_reg_internal_reg_16 : dffr port map ( Q=>LFSROUT_16, QB=>OPEN, D=>
      nx1369, CLK=>clk, R=>nx5808);
   LFSR0_reg_internal_reg_17 : dffr port map ( Q=>LFSROUT_17, QB=>OPEN, D=>
      nx1679, CLK=>clk, R=>nx5808);
   LFSR0_reg_internal_reg_18 : dffs port map ( Q=>LFSROUT_18, QB=>OPEN, D=>
      nx1669, CLK=>clk, S=>nx5808);
   LFSR0_reg_internal_reg_19 : dffr port map ( Q=>LFSROUT_19, QB=>OPEN, D=>
      nx1659, CLK=>clk, R=>nx5808);
   LFSR0_reg_internal_reg_20 : dffs port map ( Q=>LFSROUT_20, QB=>OPEN, D=>
      nx1649, CLK=>clk, S=>nx5808);
   LFSR0_reg_internal_reg_21 : dffs port map ( Q=>LFSROUT_21, QB=>OPEN, D=>
      nx1639, CLK=>clk, S=>nx5808);
   LFSR0_reg_internal_reg_22 : dffr port map ( Q=>LFSROUT_22, QB=>OPEN, D=>
      nx1629, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_23 : dffr port map ( Q=>LFSROUT_23, QB=>OPEN, D=>
      nx1619, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_24 : dffr port map ( Q=>LFSROUT_24, QB=>OPEN, D=>
      nx1609, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_25 : dffs port map ( Q=>LFSROUT_25, QB=>OPEN, D=>
      nx1599, CLK=>clk, S=>nx5806);
   LFSR0_reg_internal_reg_26 : dffr port map ( Q=>LFSROUT_26, QB=>OPEN, D=>
      nx1589, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_27 : dffr port map ( Q=>LFSROUT_27, QB=>OPEN, D=>
      nx1579, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_28 : dffs port map ( Q=>LFSROUT_28, QB=>OPEN, D=>
      nx1569, CLK=>clk, S=>nx5806);
   LFSR0_reg_internal_reg_29 : dffr port map ( Q=>LFSROUT_29, QB=>OPEN, D=>
      nx1559, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_30 : dffr port map ( Q=>LFSROUT_30, QB=>OPEN, D=>
      nx1549, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_31 : dffr port map ( Q=>LFSROUT_31, QB=>OPEN, D=>
      nx1539, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_0 : dffr port map ( Q=>LFSROUT_0, QB=>OPEN, D=>
      nx1529, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_1 : dffr port map ( Q=>LFSROUT_1, QB=>OPEN, D=>
      nx1519, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_2 : dffr port map ( Q=>LFSROUT_2, QB=>OPEN, D=>
      nx1509, CLK=>clk, R=>nx5806);
   LFSR0_reg_internal_reg_3 : dffs port map ( Q=>LFSROUT_3, QB=>OPEN, D=>
      nx1499, CLK=>clk, S=>nx5806);
   LFSR0_reg_internal_reg_4 : dffs port map ( Q=>LFSROUT_4, QB=>OPEN, D=>
      nx1489, CLK=>clk, S=>nx5806);
   LFSR0_reg_internal_reg_5 : dffs port map ( Q=>LFSROUT_5, QB=>OPEN, D=>
      nx1479, CLK=>clk, S=>nx5804);
   LFSR0_reg_internal_reg_6 : dffs port map ( Q=>LFSROUT_6, QB=>OPEN, D=>
      nx1469, CLK=>clk, S=>nx5804);
   LFSR0_reg_internal_reg_7 : dffr port map ( Q=>LFSROUT_7, QB=>OPEN, D=>
      nx1459, CLK=>clk, R=>nx5804);
   LFSR0_reg_internal_reg_8 : dffr port map ( Q=>LFSROUT_8, QB=>OPEN, D=>
      nx1449, CLK=>clk, R=>nx5804);
   LFSR0_reg_internal_reg_9 : dffs port map ( Q=>LFSROUT_9, QB=>OPEN, D=>
      nx1439, CLK=>clk, S=>nx5804);
   LFSR0_reg_internal_reg_10 : dffs port map ( Q=>LFSROUT_10, QB=>OPEN, D=>
      nx1429, CLK=>clk, S=>nx5804);
   LFSR0_reg_internal_reg_11 : dffr port map ( Q=>LFSROUT_11, QB=>OPEN, D=>
      nx1419, CLK=>clk, R=>nx5804);
   LFSR0_reg_internal_reg_12 : dffs port map ( Q=>LFSROUT_12, QB=>OPEN, D=>
      nx1409, CLK=>clk, S=>nx5804);
   LFSR0_reg_internal_reg_13 : dffr port map ( Q=>LFSROUT_13, QB=>OPEN, D=>
      nx1399, CLK=>clk, R=>nx5804);
   LFSR0_reg_internal_reg_14 : dffs port map ( Q=>LFSROUT_14, QB=>OPEN, D=>
      nx1389, CLK=>clk, S=>nx5804);
   LFSR0_reg_internal_reg_15 : dffr port map ( Q=>LFSROUT_15, QB=>OPEN, D=>
      nx1379, CLK=>clk, R=>nx5804);
   MAC0_RegMultInB_reg_Y_0 : dffr port map ( Q=>MAC0_MultB_0, QB=>OPEN, D=>
      nx698, CLK=>clk, R=>nx5808);
   ix3116 : inv01 port map ( Y=>nx3115, A=>WE);
   ix3118 : nand02 port map ( Y=>nx3117, A0=>RegOut_dup0_0, A1=>nx3115);
   MAC0_RegMultOut_reg_Y_1 : dffr port map ( Q=>MAC0_adderB_1, QB=>OPEN, D=>
      nx4000, CLK=>clk, R=>nx5808);
   ix4001 : nor02ii port map ( Y=>nx4000, A0=>nx3125, A1=>nx3137);
   ix3126 : aoi22 port map ( Y=>nx3125, A0=>nx5852, A1=>nx5848, B0=>nx5844, 
      B1=>nx5856);
   MAC0_RegMultInB_reg_Y_1 : dffr port map ( Q=>OPEN, QB=>nx3131, D=>nx672, 
      CLK=>clk, R=>nx5808);
   MAC0_RegMultInA_reg_Y_1 : dffr port map ( Q=>OPEN, QB=>nx3135, D=>nx660, 
      CLK=>clk, R=>nx5808);
   ix3144 : xnor2 port map ( Y=>nx3143, A0=>nx989, A1=>nx3145);
   ix3146 : xnor2 port map ( Y=>nx3145, A0=>MAC0_adderB_1, A1=>RegOut_dup0_1
   );
   MAC0_RegMultOut_reg_Y_2 : dffr port map ( Q=>MAC0_adderB_2, QB=>OPEN, D=>
      nx3986, CLK=>clk, R=>nx5810);
   ix3987 : aoi21 port map ( Y=>nx3986, A0=>nx3153, A1=>nx3161, B0=>nx740);
   MAC0_RegMultInA_reg_Y_2 : dffr port map ( Q=>OPEN, QB=>nx3159, D=>nx732, 
      CLK=>clk, R=>nx5808);
   ix3162 : xnor2 port map ( Y=>nx3161, A0=>nx3137, A1=>nx3163);
   ix3164 : xnor2 port map ( Y=>nx3163, A0=>nx3165, A1=>nx3167);
   ix3168 : nand02 port map ( Y=>nx3167, A0=>nx5852, A1=>nx5860);
   MAC0_RegMultInB_reg_Y_2 : dffr port map ( Q=>OPEN, QB=>nx3173, D=>nx714, 
      CLK=>clk, R=>nx5810);
   ix741 : nor03 port map ( Y=>nx740, A0=>nx3161, A1=>nx6026, A2=>nx5972);
   ix3180 : xnor2 port map ( Y=>nx3179, A0=>nx2887, A1=>nx4046);
   ix4047 : xnor2 port map ( Y=>nx4046, A0=>MAC0_adderB_2, A1=>RegOut_dup0_2
   );
   MAC0_RegMultOut_reg_Y_3 : dffr port map ( Q=>MAC0_adderB_3, QB=>OPEN, D=>
      nx3974, CLK=>clk, R=>nx5810);
   ix3975 : aoi21 port map ( Y=>nx3974, A0=>nx3189, A1=>nx3197, B0=>nx788);
   MAC0_RegMultInA_reg_Y_3 : dffr port map ( Q=>OPEN, QB=>nx3195, D=>nx780, 
      CLK=>clk, R=>nx5810);
   ix3198 : xnor2 port map ( Y=>nx3197, A0=>nx740, A1=>nx770);
   ix771 : xnor2 port map ( Y=>nx770, A0=>nx3201, A1=>nx768);
   ix769 : xnor2 port map ( Y=>nx768, A0=>nx748, A1=>nx3209);
   ix749 : aoi21 port map ( Y=>nx748, A0=>nx3167, A1=>nx3207, B0=>nx3165);
   ix3208 : nand02 port map ( Y=>nx3207, A0=>nx5852, A1=>nx5856);
   ix3210 : xnor2 port map ( Y=>nx3209, A0=>nx3211, A1=>nx3213);
   ix3214 : nand02 port map ( Y=>nx3213, A0=>nx5852, A1=>nx5868);
   MAC0_RegMultInB_reg_Y_3 : dffr port map ( Q=>OPEN, QB=>nx3219, D=>nx758, 
      CLK=>clk, R=>nx5810);
   ix789 : nor03 port map ( Y=>nx788, A0=>nx3197, A1=>nx6034, A2=>nx5972);
   ix3226 : xnor2 port map ( Y=>nx3225, A0=>nx2879, A1=>nx4062);
   ix4063 : xnor2 port map ( Y=>nx4062, A0=>MAC0_adderB_3, A1=>RegOut_dup0_3
   );
   MAC0_RegMultOut_reg_Y_4 : dffr port map ( Q=>MAC0_adderB_4, QB=>OPEN, D=>
      nx3962, CLK=>clk, R=>nx5810);
   ix3963 : aoi21 port map ( Y=>nx3962, A0=>nx3235, A1=>nx3243, B0=>nx848);
   MAC0_RegMultInA_reg_Y_4 : dffr port map ( Q=>OPEN, QB=>nx3241, D=>nx840, 
      CLK=>clk, R=>nx5810);
   ix3244 : xnor2 port map ( Y=>nx3243, A0=>nx788, A1=>nx830);
   ix831 : xnor2 port map ( Y=>nx830, A0=>nx3247, A1=>nx828);
   ix829 : xnor2 port map ( Y=>nx828, A0=>nx3251, A1=>nx826);
   ix3252 : aoi32 port map ( Y=>nx3251, A0=>nx5864, A1=>nx5848, A2=>nx768, 
      B0=>nx740, B1=>nx770);
   ix827 : xnor2 port map ( Y=>nx826, A0=>nx3255, A1=>nx824);
   ix825 : xnor2 port map ( Y=>nx824, A0=>nx804, A1=>nx3263);
   ix805 : oai32 port map ( Y=>nx804, A0=>nx6020, A1=>nx6030, A2=>nx3213, B0
      =>nx3261, B1=>nx3209);
   ix3264 : xnor2 port map ( Y=>nx3263, A0=>nx3265, A1=>nx3267);
   ix3268 : nand02 port map ( Y=>nx3267, A0=>nx5852, A1=>nx5876);
   MAC0_RegMultInB_reg_Y_4 : dffr port map ( Q=>OPEN, QB=>nx3273, D=>nx814, 
      CLK=>clk, R=>nx5810);
   ix849 : nor03 port map ( Y=>nx848, A0=>nx3243, A1=>nx6042, A2=>nx5972);
   ix3280 : xnor2 port map ( Y=>nx3279, A0=>nx2871, A1=>nx4078);
   ix4079 : xnor2 port map ( Y=>nx4078, A0=>MAC0_adderB_4, A1=>RegOut_dup0_4
   );
   MAC0_RegMultOut_reg_Y_5 : dffr port map ( Q=>MAC0_adderB_5, QB=>OPEN, D=>
      nx3950, CLK=>clk, R=>nx5810);
   ix3951 : aoi21 port map ( Y=>nx3950, A0=>nx3289, A1=>nx3297, B0=>nx920);
   MAC0_RegMultInA_reg_Y_5 : dffr port map ( Q=>OPEN, QB=>nx3295, D=>nx912, 
      CLK=>clk, R=>nx5810);
   ix3298 : xnor2 port map ( Y=>nx3297, A0=>nx848, A1=>nx902);
   ix903 : xnor2 port map ( Y=>nx902, A0=>nx3301, A1=>nx900);
   ix901 : xnor2 port map ( Y=>nx900, A0=>nx3305, A1=>nx898);
   ix3306 : aoi32 port map ( Y=>nx3305, A0=>nx5872, A1=>nx5848, A2=>nx828, 
      B0=>nx788, B1=>nx830);
   ix899 : xnor2 port map ( Y=>nx898, A0=>nx3309, A1=>nx896);
   ix897 : xnor2 port map ( Y=>nx896, A0=>nx3313, A1=>nx894);
   ix3314 : aoi32 port map ( Y=>nx3313, A0=>nx5864, A1=>nx5860, A2=>nx824, 
      B0=>nx796, B1=>nx826);
   ix895 : xnor2 port map ( Y=>nx894, A0=>nx3319, A1=>nx892);
   ix893 : xnor2 port map ( Y=>nx892, A0=>nx872, A1=>nx3331);
   ix873 : oai32 port map ( Y=>nx872, A0=>nx6020, A1=>nx6038, A2=>nx3267, B0
      =>nx3325, B1=>nx3263);
   ix3332 : xnor2 port map ( Y=>nx3331, A0=>nx3333, A1=>nx3335);
   ix3336 : nand02 port map ( Y=>nx3335, A0=>nx5852, A1=>nx5884);
   MAC0_RegMultInB_reg_Y_5 : dffr port map ( Q=>OPEN, QB=>nx3341, D=>nx882, 
      CLK=>clk, R=>nx5810);
   ix921 : nor03 port map ( Y=>nx920, A0=>nx3297, A1=>nx6050, A2=>nx5972);
   ix3348 : xnor2 port map ( Y=>nx3347, A0=>nx2863, A1=>nx4094);
   ix4095 : xnor2 port map ( Y=>nx4094, A0=>MAC0_adderB_5, A1=>RegOut_dup0_5
   );
   MAC0_RegMultOut_reg_Y_6 : dffr port map ( Q=>MAC0_adderB_6, QB=>OPEN, D=>
      nx3938, CLK=>clk, R=>nx5812);
   ix3939 : mux21 port map ( Y=>nx3938, A0=>nx3357, A1=>nx3932, S0=>nx3365);
   MAC0_RegMultInA_reg_Y_6 : dffr port map ( Q=>OPEN, QB=>nx3363, D=>nx996, 
      CLK=>clk, R=>nx5812);
   ix3366 : xnor2 port map ( Y=>nx3365, A0=>nx920, A1=>nx986);
   ix987 : xnor2 port map ( Y=>nx986, A0=>nx3369, A1=>nx984);
   ix985 : xnor2 port map ( Y=>nx984, A0=>nx3373, A1=>nx982);
   ix3374 : aoi32 port map ( Y=>nx3373, A0=>nx5880, A1=>nx5848, A2=>nx900, 
      B0=>nx848, B1=>nx902);
   ix983 : xnor2 port map ( Y=>nx982, A0=>nx3377, A1=>nx980);
   ix981 : xnor2 port map ( Y=>nx980, A0=>nx3381, A1=>nx978);
   ix3382 : aoi32 port map ( Y=>nx3381, A0=>nx5872, A1=>nx5860, A2=>nx896, 
      B0=>nx856, B1=>nx898);
   ix979 : xnor2 port map ( Y=>nx978, A0=>nx3387, A1=>nx976);
   ix977 : xnor2 port map ( Y=>nx976, A0=>nx3391, A1=>nx974);
   ix3392 : aoi32 port map ( Y=>nx3391, A0=>nx5864, A1=>nx5868, A2=>nx892, 
      B0=>nx864, B1=>nx894);
   ix975 : xnor2 port map ( Y=>nx974, A0=>nx3397, A1=>nx972);
   ix973 : xnor2 port map ( Y=>nx972, A0=>nx952, A1=>nx3409);
   ix953 : oai32 port map ( Y=>nx952, A0=>nx6020, A1=>nx6046, A2=>nx3335, B0
      =>nx3403, B1=>nx3331);
   ix3410 : xnor2 port map ( Y=>nx3409, A0=>nx3411, A1=>nx3413);
   ix3414 : nand02 port map ( Y=>nx3413, A0=>nx5852, A1=>nx5892);
   MAC0_RegMultInB_reg_Y_6 : dffr port map ( Q=>OPEN, QB=>nx3419, D=>nx962, 
      CLK=>clk, R=>nx5812);
   ix3426 : xnor2 port map ( Y=>nx3425, A0=>nx2855, A1=>nx4110);
   ix4111 : xnor2 port map ( Y=>nx4110, A0=>MAC0_adderB_6, A1=>RegOut_dup0_6
   );
   MAC0_RegMultOut_reg_Y_7 : dffr port map ( Q=>MAC0_adderB_7, QB=>OPEN, D=>
      nx3926, CLK=>clk, R=>nx5812);
   ix3927 : mux21 port map ( Y=>nx3926, A0=>nx3435, A1=>nx3920, S0=>nx3443);
   MAC0_RegMultInA_reg_Y_7 : dffr port map ( Q=>OPEN, QB=>nx3441, D=>nx1092, 
      CLK=>clk, R=>nx5812);
   ix3444 : xnor2 port map ( Y=>nx3443, A0=>nx1004, A1=>nx1082);
   ix1005 : nor03 port map ( Y=>nx1004, A0=>nx3365, A1=>nx6058, A2=>nx5972);
   ix1083 : xnor2 port map ( Y=>nx1082, A0=>nx3449, A1=>nx1080);
   ix1081 : xnor2 port map ( Y=>nx1080, A0=>nx3453, A1=>nx1078);
   ix3454 : aoi32 port map ( Y=>nx3453, A0=>nx5888, A1=>nx5848, A2=>nx984, 
      B0=>nx920, B1=>nx986);
   ix1079 : xnor2 port map ( Y=>nx1078, A0=>nx3457, A1=>nx1076);
   ix1077 : xnor2 port map ( Y=>nx1076, A0=>nx3461, A1=>nx1074);
   ix3462 : aoi32 port map ( Y=>nx3461, A0=>nx5880, A1=>nx5860, A2=>nx980, 
      B0=>nx928, B1=>nx982);
   ix1075 : xnor2 port map ( Y=>nx1074, A0=>nx3467, A1=>nx1072);
   ix1073 : xnor2 port map ( Y=>nx1072, A0=>nx3471, A1=>nx1070);
   ix3472 : aoi32 port map ( Y=>nx3471, A0=>nx5872, A1=>nx5868, A2=>nx976, 
      B0=>nx936, B1=>nx978);
   ix1071 : xnor2 port map ( Y=>nx1070, A0=>nx3477, A1=>nx1068);
   ix1069 : xnor2 port map ( Y=>nx1068, A0=>nx3481, A1=>nx1066);
   ix3482 : aoi32 port map ( Y=>nx3481, A0=>nx5864, A1=>nx5876, A2=>nx972, 
      B0=>nx944, B1=>nx974);
   ix1067 : xnor2 port map ( Y=>nx1066, A0=>nx3487, A1=>nx1064);
   ix1065 : xnor2 port map ( Y=>nx1064, A0=>nx1044, A1=>nx3499);
   ix1045 : oai32 port map ( Y=>nx1044, A0=>nx6020, A1=>nx6054, A2=>nx3413, 
      B0=>nx3493, B1=>nx3409);
   ix3500 : xnor2 port map ( Y=>nx3499, A0=>nx3501, A1=>nx3503);
   ix3504 : nand02 port map ( Y=>nx3503, A0=>nx5852, A1=>nx5900);
   MAC0_RegMultInB_reg_Y_7 : dffr port map ( Q=>OPEN, QB=>nx3509, D=>nx1054, 
      CLK=>clk, R=>nx5812);
   ix3516 : xnor2 port map ( Y=>nx3515, A0=>nx2847, A1=>nx4126);
   ix4127 : xnor2 port map ( Y=>nx4126, A0=>MAC0_adderB_7, A1=>RegOut_dup0_7
   );
   MAC0_RegMultOut_reg_Y_8 : dffr port map ( Q=>MAC0_adderB_8, QB=>OPEN, D=>
      nx3914, CLK=>clk, R=>nx5812);
   ix3915 : mux21 port map ( Y=>nx3914, A0=>nx3525, A1=>nx3908, S0=>nx3533);
   MAC0_RegMultInA_reg_Y_8 : dffr port map ( Q=>OPEN, QB=>nx3531, D=>nx1200, 
      CLK=>clk, R=>nx5812);
   ix3534 : xnor2 port map ( Y=>nx3533, A0=>nx1100, A1=>nx1190);
   ix1101 : nor03 port map ( Y=>nx1100, A0=>nx3443, A1=>nx6066, A2=>nx5972);
   ix1191 : xnor2 port map ( Y=>nx1190, A0=>nx3539, A1=>nx1188);
   ix1189 : xnor2 port map ( Y=>nx1188, A0=>nx3543, A1=>nx1186);
   ix3544 : aoi32 port map ( Y=>nx3543, A0=>nx5896, A1=>nx5848, A2=>nx1080, 
      B0=>nx1004, B1=>nx1082);
   ix1187 : xnor2 port map ( Y=>nx1186, A0=>nx3547, A1=>nx1184);
   ix1185 : xnor2 port map ( Y=>nx1184, A0=>nx3551, A1=>nx1182);
   ix3552 : aoi32 port map ( Y=>nx3551, A0=>nx5888, A1=>nx5860, A2=>nx1076, 
      B0=>nx1012, B1=>nx1078);
   ix1183 : xnor2 port map ( Y=>nx1182, A0=>nx3557, A1=>nx1180);
   ix1181 : xnor2 port map ( Y=>nx1180, A0=>nx3561, A1=>nx1178);
   ix3562 : aoi32 port map ( Y=>nx3561, A0=>nx5880, A1=>nx5868, A2=>nx1072, 
      B0=>nx1020, B1=>nx1074);
   ix1179 : xnor2 port map ( Y=>nx1178, A0=>nx3567, A1=>nx1176);
   ix1177 : xnor2 port map ( Y=>nx1176, A0=>nx3571, A1=>nx1174);
   ix3572 : aoi32 port map ( Y=>nx3571, A0=>nx5872, A1=>nx5876, A2=>nx1068, 
      B0=>nx1028, B1=>nx1070);
   ix1175 : xnor2 port map ( Y=>nx1174, A0=>nx3577, A1=>nx1172);
   ix1173 : xnor2 port map ( Y=>nx1172, A0=>nx3581, A1=>nx1170);
   ix3582 : aoi32 port map ( Y=>nx3581, A0=>nx5864, A1=>nx5884, A2=>nx1064, 
      B0=>nx1036, B1=>nx1066);
   ix1171 : xnor2 port map ( Y=>nx1170, A0=>nx3587, A1=>nx1168);
   ix1169 : xnor2 port map ( Y=>nx1168, A0=>nx1148, A1=>nx3599);
   ix1149 : oai32 port map ( Y=>nx1148, A0=>nx6020, A1=>nx6062, A2=>nx3503, 
      B0=>nx3593, B1=>nx3499);
   ix3600 : xnor2 port map ( Y=>nx3599, A0=>nx3601, A1=>nx3603);
   ix3604 : nand02 port map ( Y=>nx3603, A0=>nx5852, A1=>nx5908);
   MAC0_RegMultInB_reg_Y_8 : dffr port map ( Q=>OPEN, QB=>nx3609, D=>nx1158, 
      CLK=>clk, R=>nx5812);
   ix3616 : xnor2 port map ( Y=>nx3615, A0=>nx2839, A1=>nx4142);
   ix4143 : xnor2 port map ( Y=>nx4142, A0=>MAC0_adderB_8, A1=>RegOut_dup0_8
   );
   MAC0_RegMultOut_reg_Y_9 : dffr port map ( Q=>MAC0_adderB_9, QB=>OPEN, D=>
      nx3902, CLK=>clk, R=>nx5812);
   ix3903 : mux21 port map ( Y=>nx3902, A0=>nx3625, A1=>nx3896, S0=>nx3633);
   MAC0_RegMultInA_reg_Y_9 : dffr port map ( Q=>OPEN, QB=>nx3631, D=>nx1320, 
      CLK=>clk, R=>nx5812);
   ix3634 : xnor2 port map ( Y=>nx3633, A0=>nx1208, A1=>nx1310);
   ix1209 : nor03 port map ( Y=>nx1208, A0=>nx3533, A1=>nx6074, A2=>nx5972);
   ix1311 : xnor2 port map ( Y=>nx1310, A0=>nx3639, A1=>nx1308);
   ix1309 : xnor2 port map ( Y=>nx1308, A0=>nx3643, A1=>nx1306);
   ix3644 : aoi32 port map ( Y=>nx3643, A0=>nx5904, A1=>nx5850, A2=>nx1188, 
      B0=>nx1100, B1=>nx1190);
   ix1307 : xnor2 port map ( Y=>nx1306, A0=>nx3647, A1=>nx1304);
   ix1305 : xnor2 port map ( Y=>nx1304, A0=>nx3651, A1=>nx1302);
   ix3652 : aoi32 port map ( Y=>nx3651, A0=>nx5896, A1=>nx5860, A2=>nx1184, 
      B0=>nx1108, B1=>nx1186);
   ix1303 : xnor2 port map ( Y=>nx1302, A0=>nx3657, A1=>nx1300);
   ix1301 : xnor2 port map ( Y=>nx1300, A0=>nx3661, A1=>nx1298);
   ix3662 : aoi32 port map ( Y=>nx3661, A0=>nx5888, A1=>nx5868, A2=>nx1180, 
      B0=>nx1116, B1=>nx1182);
   ix1299 : xnor2 port map ( Y=>nx1298, A0=>nx3667, A1=>nx1296);
   ix1297 : xnor2 port map ( Y=>nx1296, A0=>nx3671, A1=>nx1294);
   ix3672 : aoi32 port map ( Y=>nx3671, A0=>nx5880, A1=>nx5876, A2=>nx1176, 
      B0=>nx1124, B1=>nx1178);
   ix1295 : xnor2 port map ( Y=>nx1294, A0=>nx3677, A1=>nx1292);
   ix1293 : xnor2 port map ( Y=>nx1292, A0=>nx3681, A1=>nx1290);
   ix3682 : aoi32 port map ( Y=>nx3681, A0=>nx5872, A1=>nx5884, A2=>nx1172, 
      B0=>nx1132, B1=>nx1174);
   ix1291 : xnor2 port map ( Y=>nx1290, A0=>nx3687, A1=>nx1288);
   ix1289 : xnor2 port map ( Y=>nx1288, A0=>nx3691, A1=>nx1286);
   ix3692 : aoi32 port map ( Y=>nx3691, A0=>nx5864, A1=>nx5892, A2=>nx1168, 
      B0=>nx1140, B1=>nx1170);
   ix1287 : xnor2 port map ( Y=>nx1286, A0=>nx3697, A1=>nx1284);
   ix1285 : xnor2 port map ( Y=>nx1284, A0=>nx1264, A1=>nx3709);
   ix1265 : oai32 port map ( Y=>nx1264, A0=>nx6020, A1=>nx6070, A2=>nx3603, 
      B0=>nx3703, B1=>nx3599);
   ix3710 : xnor2 port map ( Y=>nx3709, A0=>nx3711, A1=>nx3713);
   ix3714 : nand02 port map ( Y=>nx3713, A0=>nx5852, A1=>nx5916);
   MAC0_RegMultInB_reg_Y_9 : dffr port map ( Q=>OPEN, QB=>nx3719, D=>nx1274, 
      CLK=>clk, R=>nx5812);
   ix3726 : xnor2 port map ( Y=>nx3725, A0=>nx2831, A1=>nx4158);
   ix4159 : xnor2 port map ( Y=>nx4158, A0=>MAC0_adderB_9, A1=>RegOut_dup0_9
   );
   MAC0_RegMultOut_reg_Y_10 : dffr port map ( Q=>MAC0_adderB_10, QB=>OPEN, D
      =>nx3890, CLK=>clk, R=>nx5814);
   ix3891 : mux21 port map ( Y=>nx3890, A0=>nx3735, A1=>nx3884, S0=>nx3743);
   MAC0_RegMultInA_reg_Y_10 : dffr port map ( Q=>OPEN, QB=>nx3741, D=>nx1452, 
      CLK=>clk, R=>nx5814);
   ix3744 : xnor2 port map ( Y=>nx3743, A0=>nx1328, A1=>nx1442);
   ix1329 : nor03 port map ( Y=>nx1328, A0=>nx3633, A1=>nx6082, A2=>nx5972);
   ix1443 : xnor2 port map ( Y=>nx1442, A0=>nx3749, A1=>nx1440);
   ix1441 : xnor2 port map ( Y=>nx1440, A0=>nx3753, A1=>nx1438);
   ix3754 : aoi32 port map ( Y=>nx3753, A0=>nx5912, A1=>nx5850, A2=>nx1308, 
      B0=>nx1208, B1=>nx1310);
   ix1439 : xnor2 port map ( Y=>nx1438, A0=>nx3756, A1=>nx1436);
   ix1437 : xnor2 port map ( Y=>nx1436, A0=>nx3759, A1=>nx1434);
   ix3760 : aoi32 port map ( Y=>nx3759, A0=>nx5904, A1=>nx5860, A2=>nx1304, 
      B0=>nx1216, B1=>nx1306);
   ix1435 : xnor2 port map ( Y=>nx1434, A0=>nx3763, A1=>nx1432);
   ix1433 : xnor2 port map ( Y=>nx1432, A0=>nx3767, A1=>nx1430);
   ix3768 : aoi32 port map ( Y=>nx3767, A0=>nx5896, A1=>nx5868, A2=>nx1300, 
      B0=>nx1224, B1=>nx1302);
   ix1431 : xnor2 port map ( Y=>nx1430, A0=>nx3771, A1=>nx1428);
   ix1429 : xnor2 port map ( Y=>nx1428, A0=>nx3774, A1=>nx1426);
   ix3775 : aoi32 port map ( Y=>nx3774, A0=>nx5888, A1=>nx5876, A2=>nx1296, 
      B0=>nx1232, B1=>nx1298);
   ix1427 : xnor2 port map ( Y=>nx1426, A0=>nx3779, A1=>nx1424);
   ix1425 : xnor2 port map ( Y=>nx1424, A0=>nx3783, A1=>nx1422);
   ix3784 : aoi32 port map ( Y=>nx3783, A0=>nx5880, A1=>nx5884, A2=>nx1292, 
      B0=>nx1240, B1=>nx1294);
   ix1423 : xnor2 port map ( Y=>nx1422, A0=>nx3787, A1=>nx1420);
   ix1421 : xnor2 port map ( Y=>nx1420, A0=>nx3791, A1=>nx1418);
   ix3792 : aoi32 port map ( Y=>nx3791, A0=>nx5872, A1=>nx5892, A2=>nx1288, 
      B0=>nx1248, B1=>nx1290);
   ix1419 : xnor2 port map ( Y=>nx1418, A0=>nx3795, A1=>nx1416);
   ix1417 : xnor2 port map ( Y=>nx1416, A0=>nx3798, A1=>nx1414);
   ix3799 : aoi32 port map ( Y=>nx3798, A0=>nx5864, A1=>nx5900, A2=>nx1284, 
      B0=>nx1256, B1=>nx1286);
   ix1415 : xnor2 port map ( Y=>nx1414, A0=>nx3803, A1=>nx1412);
   ix1413 : xnor2 port map ( Y=>nx1412, A0=>nx1392, A1=>nx3811);
   ix1393 : oai32 port map ( Y=>nx1392, A0=>nx6020, A1=>nx6078, A2=>nx3713, 
      B0=>nx3807, B1=>nx3709);
   ix3812 : xnor2 port map ( Y=>nx3811, A0=>nx3813, A1=>nx3815);
   ix3816 : nand02 port map ( Y=>nx3815, A0=>nx5852, A1=>nx5924);
   MAC0_RegMultInB_reg_Y_10 : dffr port map ( Q=>OPEN, QB=>nx3819, D=>nx1402, 
      CLK=>clk, R=>nx5814);
   ix3824 : xnor2 port map ( Y=>nx3823, A0=>nx2823, A1=>nx4174);
   ix4175 : xnor2 port map ( Y=>nx4174, A0=>MAC0_adderB_10, A1=>
      RegOut_dup0_10);
   MAC0_RegMultOut_reg_Y_11 : dffr port map ( Q=>MAC0_adderB_11, QB=>OPEN, D
      =>nx3878, CLK=>clk, R=>nx5814);
   ix3879 : mux21 port map ( Y=>nx3878, A0=>nx3833, A1=>nx3872, S0=>nx3839);
   MAC0_RegMultInA_reg_Y_11 : dffr port map ( Q=>OPEN, QB=>nx3837, D=>nx1596, 
      CLK=>clk, R=>nx5814);
   ix3840 : xnor2 port map ( Y=>nx3839, A0=>nx1460, A1=>nx1586);
   ix1461 : nor03 port map ( Y=>nx1460, A0=>nx3743, A1=>nx6090, A2=>nx5972);
   ix1587 : xnor2 port map ( Y=>nx1586, A0=>nx3845, A1=>nx1584);
   ix1585 : xnor2 port map ( Y=>nx1584, A0=>nx3849, A1=>nx1582);
   ix3850 : aoi32 port map ( Y=>nx3849, A0=>nx5920, A1=>nx5850, A2=>nx1440, 
      B0=>nx1328, B1=>nx1442);
   ix1583 : xnor2 port map ( Y=>nx1582, A0=>nx3853, A1=>nx1580);
   ix1581 : xnor2 port map ( Y=>nx1580, A0=>nx3857, A1=>nx1578);
   ix3858 : aoi32 port map ( Y=>nx3857, A0=>nx5912, A1=>nx5862, A2=>nx1436, 
      B0=>nx1336, B1=>nx1438);
   ix1579 : xnor2 port map ( Y=>nx1578, A0=>nx3861, A1=>nx1576);
   ix1577 : xnor2 port map ( Y=>nx1576, A0=>nx3865, A1=>nx1574);
   ix3866 : aoi32 port map ( Y=>nx3865, A0=>nx5904, A1=>nx5868, A2=>nx1432, 
      B0=>nx1344, B1=>nx1434);
   ix1575 : xnor2 port map ( Y=>nx1574, A0=>nx3870, A1=>nx1572);
   ix1573 : xnor2 port map ( Y=>nx1572, A0=>nx3873, A1=>nx1570);
   ix3874 : aoi32 port map ( Y=>nx3873, A0=>nx5896, A1=>nx5876, A2=>nx1428, 
      B0=>nx1352, B1=>nx1430);
   ix1571 : xnor2 port map ( Y=>nx1570, A0=>nx3879, A1=>nx1568);
   ix1569 : xnor2 port map ( Y=>nx1568, A0=>nx3882, A1=>nx1566);
   ix3883 : aoi32 port map ( Y=>nx3882, A0=>nx5888, A1=>nx5884, A2=>nx1424, 
      B0=>nx1360, B1=>nx1426);
   ix1567 : xnor2 port map ( Y=>nx1566, A0=>nx3887, A1=>nx1564);
   ix1565 : xnor2 port map ( Y=>nx1564, A0=>nx3891, A1=>nx1562);
   ix3892 : aoi32 port map ( Y=>nx3891, A0=>nx5880, A1=>nx5892, A2=>nx1420, 
      B0=>nx1368, B1=>nx1422);
   ix1563 : xnor2 port map ( Y=>nx1562, A0=>nx3895, A1=>nx1560);
   ix1561 : xnor2 port map ( Y=>nx1560, A0=>nx3899, A1=>nx1558);
   ix3900 : aoi32 port map ( Y=>nx3899, A0=>nx5872, A1=>nx5900, A2=>nx1416, 
      B0=>nx1376, B1=>nx1418);
   ix1559 : xnor2 port map ( Y=>nx1558, A0=>nx3905, A1=>nx1556);
   ix1557 : xnor2 port map ( Y=>nx1556, A0=>nx3909, A1=>nx1554);
   ix3910 : aoi32 port map ( Y=>nx3909, A0=>nx5866, A1=>nx5908, A2=>nx1412, 
      B0=>nx1384, B1=>nx1414);
   ix1555 : xnor2 port map ( Y=>nx1554, A0=>nx3915, A1=>nx1552);
   ix1553 : xnor2 port map ( Y=>nx1552, A0=>nx1532, A1=>nx3925);
   ix1533 : oai32 port map ( Y=>nx1532, A0=>nx6020, A1=>nx6086, A2=>nx3815, 
      B0=>nx3919, B1=>nx3811);
   ix3926 : xnor2 port map ( Y=>nx3925, A0=>nx3927, A1=>nx3929);
   ix3930 : nand02 port map ( Y=>nx3929, A0=>nx5852, A1=>nx5932);
   MAC0_RegMultInB_reg_Y_11 : dffr port map ( Q=>OPEN, QB=>nx3933, D=>nx1542, 
      CLK=>clk, R=>nx5814);
   ix3940 : xnor2 port map ( Y=>nx3939, A0=>nx2815, A1=>nx4190);
   ix4191 : xnor2 port map ( Y=>nx4190, A0=>MAC0_adderB_11, A1=>
      RegOut_dup0_11);
   MAC0_RegMultOut_reg_Y_12 : dffr port map ( Q=>MAC0_adderB_12, QB=>OPEN, D
      =>nx3866, CLK=>clk, R=>nx5814);
   ix3867 : mux21 port map ( Y=>nx3866, A0=>nx3947, A1=>nx3860, S0=>nx3955);
   MAC0_RegMultInA_reg_Y_12 : dffr port map ( Q=>OPEN, QB=>nx3953, D=>nx1752, 
      CLK=>clk, R=>nx5814);
   ix3956 : xnor2 port map ( Y=>nx3955, A0=>nx1604, A1=>nx1742);
   ix1605 : nor03 port map ( Y=>nx1604, A0=>nx3839, A1=>nx6098, A2=>nx6140);
   ix1743 : xnor2 port map ( Y=>nx1742, A0=>nx3961, A1=>nx1740);
   ix1741 : xnor2 port map ( Y=>nx1740, A0=>nx3965, A1=>nx1738);
   ix3966 : aoi32 port map ( Y=>nx3965, A0=>nx5928, A1=>nx5850, A2=>nx1584, 
      B0=>nx1460, B1=>nx1586);
   ix1739 : xnor2 port map ( Y=>nx1738, A0=>nx3969, A1=>nx1736);
   ix1737 : xnor2 port map ( Y=>nx1736, A0=>nx3973, A1=>nx1734);
   ix3974 : aoi32 port map ( Y=>nx3973, A0=>nx5920, A1=>nx5862, A2=>nx1580, 
      B0=>nx1468, B1=>nx1582);
   ix1735 : xnor2 port map ( Y=>nx1734, A0=>nx3978, A1=>nx1732);
   ix1733 : xnor2 port map ( Y=>nx1732, A0=>nx3981, A1=>nx1730);
   ix3982 : aoi32 port map ( Y=>nx3981, A0=>nx5912, A1=>nx5870, A2=>nx1576, 
      B0=>nx1476, B1=>nx1578);
   ix1731 : xnor2 port map ( Y=>nx1730, A0=>nx3987, A1=>nx1728);
   ix1729 : xnor2 port map ( Y=>nx1728, A0=>nx3990, A1=>nx1726);
   ix3991 : aoi32 port map ( Y=>nx3990, A0=>nx5904, A1=>nx5876, A2=>nx1572, 
      B0=>nx1484, B1=>nx1574);
   ix1727 : xnor2 port map ( Y=>nx1726, A0=>nx3995, A1=>nx1724);
   ix1725 : xnor2 port map ( Y=>nx1724, A0=>nx3999, A1=>nx1722);
   ix4000 : aoi32 port map ( Y=>nx3999, A0=>nx5896, A1=>nx5884, A2=>nx1568, 
      B0=>nx1492, B1=>nx1570);
   ix1723 : xnor2 port map ( Y=>nx1722, A0=>nx4004, A1=>nx1720);
   ix1721 : xnor2 port map ( Y=>nx1720, A0=>nx4007, A1=>nx1718);
   ix4008 : aoi32 port map ( Y=>nx4007, A0=>nx5888, A1=>nx5892, A2=>nx1564, 
      B0=>nx1500, B1=>nx1566);
   ix1719 : xnor2 port map ( Y=>nx1718, A0=>nx4011, A1=>nx1716);
   ix1717 : xnor2 port map ( Y=>nx1716, A0=>nx4015, A1=>nx1714);
   ix4016 : aoi32 port map ( Y=>nx4015, A0=>nx5880, A1=>nx5900, A2=>nx1560, 
      B0=>nx1508, B1=>nx1562);
   ix1715 : xnor2 port map ( Y=>nx1714, A0=>nx4019, A1=>nx1712);
   ix1713 : xnor2 port map ( Y=>nx1712, A0=>nx4023, A1=>nx1710);
   ix4024 : aoi32 port map ( Y=>nx4023, A0=>nx5874, A1=>nx5908, A2=>nx1556, 
      B0=>nx1516, B1=>nx1558);
   ix1711 : xnor2 port map ( Y=>nx1710, A0=>nx4027, A1=>nx1708);
   ix1709 : xnor2 port map ( Y=>nx1708, A0=>nx4031, A1=>nx1706);
   ix4032 : aoi32 port map ( Y=>nx4031, A0=>nx5866, A1=>nx5916, A2=>nx1552, 
      B0=>nx1524, B1=>nx1554);
   ix1707 : xnor2 port map ( Y=>nx1706, A0=>nx4037, A1=>nx1704);
   ix1705 : xnor2 port map ( Y=>nx1704, A0=>nx1684, A1=>nx4047);
   ix1685 : oai32 port map ( Y=>nx1684, A0=>nx6020, A1=>nx6094, A2=>nx3929, 
      B0=>nx4043, B1=>nx3925);
   ix4048 : xnor2 port map ( Y=>nx4047, A0=>nx4049, A1=>nx4051);
   ix4052 : nand02 port map ( Y=>nx4051, A0=>nx5852, A1=>nx5940);
   MAC0_RegMultInB_reg_Y_12 : dffr port map ( Q=>OPEN, QB=>nx4057, D=>nx1694, 
      CLK=>clk, R=>nx5814);
   ix4062 : xnor2 port map ( Y=>nx4061, A0=>nx2807, A1=>nx4206);
   ix4207 : xnor2 port map ( Y=>nx4206, A0=>MAC0_adderB_12, A1=>
      RegOut_dup0_12);
   MAC0_RegMultOut_reg_Y_13 : dffr port map ( Q=>MAC0_adderB_13, QB=>OPEN, D
      =>nx3854, CLK=>clk, R=>nx5816);
   ix3855 : mux21 port map ( Y=>nx3854, A0=>nx4071, A1=>nx3848, S0=>nx4079);
   MAC0_RegMultInA_reg_Y_13 : dffr port map ( Q=>OPEN, QB=>nx4076, D=>nx1920, 
      CLK=>clk, R=>nx5814);
   ix4080 : xnor2 port map ( Y=>nx4079, A0=>nx1760, A1=>nx1910);
   ix1761 : nor03 port map ( Y=>nx1760, A0=>nx3955, A1=>nx6106, A2=>nx6140);
   ix1911 : xnor2 port map ( Y=>nx1910, A0=>nx4085, A1=>nx1908);
   ix1909 : xnor2 port map ( Y=>nx1908, A0=>nx4089, A1=>nx1906);
   ix4090 : aoi32 port map ( Y=>nx4089, A0=>nx5936, A1=>nx5850, A2=>nx1740, 
      B0=>nx1604, B1=>nx1742);
   ix1907 : xnor2 port map ( Y=>nx1906, A0=>nx4092, A1=>nx1904);
   ix1905 : xnor2 port map ( Y=>nx1904, A0=>nx4095, A1=>nx1902);
   ix4096 : aoi32 port map ( Y=>nx4095, A0=>nx5928, A1=>nx5862, A2=>nx1736, 
      B0=>nx1612, B1=>nx1738);
   ix1903 : xnor2 port map ( Y=>nx1902, A0=>nx4101, A1=>nx1900);
   ix1901 : xnor2 port map ( Y=>nx1900, A0=>nx4105, A1=>nx1898);
   ix4106 : aoi32 port map ( Y=>nx4105, A0=>nx5920, A1=>nx5870, A2=>nx1732, 
      B0=>nx1620, B1=>nx1734);
   ix1899 : xnor2 port map ( Y=>nx1898, A0=>nx4109, A1=>nx1896);
   ix1897 : xnor2 port map ( Y=>nx1896, A0=>nx4113, A1=>nx1894);
   ix4114 : aoi32 port map ( Y=>nx4113, A0=>nx5912, A1=>nx5878, A2=>nx1728, 
      B0=>nx1628, B1=>nx1730);
   ix1895 : xnor2 port map ( Y=>nx1894, A0=>nx4119, A1=>nx1892);
   ix1893 : xnor2 port map ( Y=>nx1892, A0=>nx4123, A1=>nx1890);
   ix4124 : aoi32 port map ( Y=>nx4123, A0=>nx5904, A1=>nx5884, A2=>nx1724, 
      B0=>nx1636, B1=>nx1726);
   ix1891 : xnor2 port map ( Y=>nx1890, A0=>nx4127, A1=>nx1888);
   ix1889 : xnor2 port map ( Y=>nx1888, A0=>nx4131, A1=>nx1886);
   ix4132 : aoi32 port map ( Y=>nx4131, A0=>nx5896, A1=>nx5892, A2=>nx1720, 
      B0=>nx1644, B1=>nx1722);
   ix1887 : xnor2 port map ( Y=>nx1886, A0=>nx4137, A1=>nx1884);
   ix1885 : xnor2 port map ( Y=>nx1884, A0=>nx4140, A1=>nx1882);
   ix4141 : aoi32 port map ( Y=>nx4140, A0=>nx5888, A1=>nx5900, A2=>nx1716, 
      B0=>nx1652, B1=>nx1718);
   ix1883 : xnor2 port map ( Y=>nx1882, A0=>nx4145, A1=>nx1880);
   ix1881 : xnor2 port map ( Y=>nx1880, A0=>nx4149, A1=>nx1878);
   ix4150 : aoi32 port map ( Y=>nx4149, A0=>nx5882, A1=>nx5908, A2=>nx1712, 
      B0=>nx1660, B1=>nx1714);
   ix1879 : xnor2 port map ( Y=>nx1878, A0=>nx4155, A1=>nx1876);
   ix1877 : xnor2 port map ( Y=>nx1876, A0=>nx4159, A1=>nx1874);
   ix4160 : aoi32 port map ( Y=>nx4159, A0=>nx5874, A1=>nx5916, A2=>nx1708, 
      B0=>nx1668, B1=>nx1710);
   ix1875 : xnor2 port map ( Y=>nx1874, A0=>nx4165, A1=>nx1872);
   ix1873 : xnor2 port map ( Y=>nx1872, A0=>nx4169, A1=>nx1870);
   ix4170 : aoi32 port map ( Y=>nx4169, A0=>nx5866, A1=>nx5924, A2=>nx1704, 
      B0=>nx1676, B1=>nx1706);
   ix1871 : xnor2 port map ( Y=>nx1870, A0=>nx4173, A1=>nx1868);
   ix1869 : xnor2 port map ( Y=>nx1868, A0=>nx1848, A1=>nx4185);
   ix1849 : oai32 port map ( Y=>nx1848, A0=>nx6020, A1=>nx6102, A2=>nx4051, 
      B0=>nx4179, B1=>nx4047);
   ix4186 : xnor2 port map ( Y=>nx4185, A0=>nx4187, A1=>nx4189);
   ix4190 : nand02 port map ( Y=>nx4189, A0=>nx5852, A1=>nx5948);
   MAC0_RegMultInB_reg_Y_13 : dffr port map ( Q=>OPEN, QB=>nx4195, D=>nx1858, 
      CLK=>clk, R=>nx5814);
   ix4202 : xnor2 port map ( Y=>nx4201, A0=>nx2799, A1=>nx4222);
   ix4223 : xnor2 port map ( Y=>nx4222, A0=>MAC0_adderB_13, A1=>
      RegOut_dup0_13);
   MAC0_RegMultOut_reg_Y_14 : dffr port map ( Q=>MAC0_adderB_14, QB=>OPEN, D
      =>nx3842, CLK=>clk, R=>nx5816);
   ix3843 : mux21 port map ( Y=>nx3842, A0=>nx4209, A1=>nx3836, S0=>nx4217);
   MAC0_RegMultInA_reg_Y_14 : dffr port map ( Q=>OPEN, QB=>nx4215, D=>nx2100, 
      CLK=>clk, R=>nx5816);
   ix4218 : xnor2 port map ( Y=>nx4217, A0=>nx1928, A1=>nx2090);
   ix1929 : nor03 port map ( Y=>nx1928, A0=>nx4079, A1=>nx6114, A2=>nx6140);
   ix2091 : xnor2 port map ( Y=>nx2090, A0=>nx4221, A1=>nx2088);
   ix2089 : xnor2 port map ( Y=>nx2088, A0=>nx4225, A1=>nx2086);
   ix4226 : aoi32 port map ( Y=>nx4225, A0=>nx5944, A1=>nx5850, A2=>nx1908, 
      B0=>nx1760, B1=>nx1910);
   ix2087 : xnor2 port map ( Y=>nx2086, A0=>nx4229, A1=>nx2084);
   ix2085 : xnor2 port map ( Y=>nx2084, A0=>nx4233, A1=>nx2082);
   ix4234 : aoi32 port map ( Y=>nx4233, A0=>nx5936, A1=>nx5862, A2=>nx1904, 
      B0=>nx1768, B1=>nx1906);
   ix2083 : xnor2 port map ( Y=>nx2082, A0=>nx4237, A1=>nx2080);
   ix2081 : xnor2 port map ( Y=>nx2080, A0=>nx4241, A1=>nx2078);
   ix4242 : aoi32 port map ( Y=>nx4241, A0=>nx5928, A1=>nx5870, A2=>nx1900, 
      B0=>nx1776, B1=>nx1902);
   ix2079 : xnor2 port map ( Y=>nx2078, A0=>nx4247, A1=>nx2076);
   ix2077 : xnor2 port map ( Y=>nx2076, A0=>nx4251, A1=>nx2074);
   ix4252 : aoi32 port map ( Y=>nx4251, A0=>nx5920, A1=>nx5878, A2=>nx1896, 
      B0=>nx1784, B1=>nx1898);
   ix2075 : xnor2 port map ( Y=>nx2074, A0=>nx4255, A1=>nx2072);
   ix2073 : xnor2 port map ( Y=>nx2072, A0=>nx4259, A1=>nx2070);
   ix4260 : aoi32 port map ( Y=>nx4259, A0=>nx5912, A1=>nx5886, A2=>nx1892, 
      B0=>nx1792, B1=>nx1894);
   ix2071 : xnor2 port map ( Y=>nx2070, A0=>nx4265, A1=>nx2068);
   ix2069 : xnor2 port map ( Y=>nx2068, A0=>nx4268, A1=>nx2066);
   ix4269 : aoi32 port map ( Y=>nx4268, A0=>nx5904, A1=>nx5892, A2=>nx1888, 
      B0=>nx1800, B1=>nx1890);
   ix2067 : xnor2 port map ( Y=>nx2066, A0=>nx4273, A1=>nx2064);
   ix2065 : xnor2 port map ( Y=>nx2064, A0=>nx4277, A1=>nx2062);
   ix4278 : aoi32 port map ( Y=>nx4277, A0=>nx5896, A1=>nx5900, A2=>nx1884, 
      B0=>nx1808, B1=>nx1886);
   ix2063 : xnor2 port map ( Y=>nx2062, A0=>nx4283, A1=>nx2060);
   ix2061 : xnor2 port map ( Y=>nx2060, A0=>nx4287, A1=>nx2058);
   ix4288 : aoi32 port map ( Y=>nx4287, A0=>nx5890, A1=>nx5908, A2=>nx1880, 
      B0=>nx1816, B1=>nx1882);
   ix2059 : xnor2 port map ( Y=>nx2058, A0=>nx4293, A1=>nx2056);
   ix2057 : xnor2 port map ( Y=>nx2056, A0=>nx4297, A1=>nx2054);
   ix4298 : aoi32 port map ( Y=>nx4297, A0=>nx5882, A1=>nx5916, A2=>nx1876, 
      B0=>nx1824, B1=>nx1878);
   ix2055 : xnor2 port map ( Y=>nx2054, A0=>nx4301, A1=>nx2052);
   ix2053 : xnor2 port map ( Y=>nx2052, A0=>nx4305, A1=>nx2050);
   ix4306 : aoi32 port map ( Y=>nx4305, A0=>nx5874, A1=>nx5924, A2=>nx1872, 
      B0=>nx1832, B1=>nx1874);
   ix2051 : xnor2 port map ( Y=>nx2050, A0=>nx4311, A1=>nx2048);
   ix2049 : xnor2 port map ( Y=>nx2048, A0=>nx4315, A1=>nx2046);
   ix4316 : aoi32 port map ( Y=>nx4315, A0=>nx5866, A1=>nx5932, A2=>nx1868, 
      B0=>nx1840, B1=>nx1870);
   ix2047 : xnor2 port map ( Y=>nx2046, A0=>nx4319, A1=>nx2044);
   ix2045 : xnor2 port map ( Y=>nx2044, A0=>nx2024, A1=>nx4331);
   ix2025 : oai32 port map ( Y=>nx2024, A0=>nx6020, A1=>nx6110, A2=>nx4189, 
      B0=>nx4325, B1=>nx4185);
   ix4332 : xnor2 port map ( Y=>nx4331, A0=>nx4333, A1=>nx4335);
   ix4336 : nand02 port map ( Y=>nx4335, A0=>nx5854, A1=>nx5956);
   MAC0_RegMultInB_reg_Y_14 : dffr port map ( Q=>OPEN, QB=>nx4341, D=>nx2034, 
      CLK=>clk, R=>nx5816);
   ix4348 : xnor2 port map ( Y=>nx4347, A0=>nx2791, A1=>nx4238);
   ix4239 : xnor2 port map ( Y=>nx4238, A0=>MAC0_adderB_14, A1=>
      RegOut_dup0_14);
   MAC0_RegMultOut_reg_Y_15 : dffr port map ( Q=>MAC0_adderB_15, QB=>OPEN, D
      =>nx3830, CLK=>clk, R=>nx5816);
   ix3831 : mux21 port map ( Y=>nx3830, A0=>nx4357, A1=>nx3824, S0=>nx4365);
   MAC0_RegMultInA_reg_Y_15 : dffr port map ( Q=>OPEN, QB=>nx4363, D=>nx2292, 
      CLK=>clk, R=>nx5816);
   ix4366 : xnor2 port map ( Y=>nx4365, A0=>nx2108, A1=>nx2282);
   ix2109 : nor03 port map ( Y=>nx2108, A0=>nx4217, A1=>nx6122, A2=>nx6140);
   ix2283 : xnor2 port map ( Y=>nx2282, A0=>nx4371, A1=>nx2280);
   ix2281 : xnor2 port map ( Y=>nx2280, A0=>nx4375, A1=>nx2278);
   ix4376 : aoi32 port map ( Y=>nx4375, A0=>nx5952, A1=>nx5850, A2=>nx2088, 
      B0=>nx1928, B1=>nx2090);
   ix2279 : xnor2 port map ( Y=>nx2278, A0=>nx4379, A1=>nx2276);
   ix2277 : xnor2 port map ( Y=>nx2276, A0=>nx4383, A1=>nx2274);
   ix4384 : aoi32 port map ( Y=>nx4383, A0=>nx5944, A1=>nx5862, A2=>nx2084, 
      B0=>nx1936, B1=>nx2086);
   ix2275 : xnor2 port map ( Y=>nx2274, A0=>nx4389, A1=>nx2272);
   ix2273 : xnor2 port map ( Y=>nx2272, A0=>nx4393, A1=>nx2270);
   ix4394 : aoi32 port map ( Y=>nx4393, A0=>nx5936, A1=>nx5870, A2=>nx2080, 
      B0=>nx1944, B1=>nx2082);
   ix2271 : xnor2 port map ( Y=>nx2270, A0=>nx4397, A1=>nx2268);
   ix2269 : xnor2 port map ( Y=>nx2268, A0=>nx4401, A1=>nx2266);
   ix4402 : aoi32 port map ( Y=>nx4401, A0=>nx5928, A1=>nx5878, A2=>nx2076, 
      B0=>nx1952, B1=>nx2078);
   ix2267 : xnor2 port map ( Y=>nx2266, A0=>nx4407, A1=>nx2264);
   ix2265 : xnor2 port map ( Y=>nx2264, A0=>nx4411, A1=>nx2262);
   ix4412 : aoi32 port map ( Y=>nx4411, A0=>nx5920, A1=>nx5886, A2=>nx2072, 
      B0=>nx1960, B1=>nx2074);
   ix2263 : xnor2 port map ( Y=>nx2262, A0=>nx4415, A1=>nx2260);
   ix2261 : xnor2 port map ( Y=>nx2260, A0=>nx4419, A1=>nx2258);
   ix4420 : aoi32 port map ( Y=>nx4419, A0=>nx5912, A1=>nx5894, A2=>nx2068, 
      B0=>nx1968, B1=>nx2070);
   ix2259 : xnor2 port map ( Y=>nx2258, A0=>nx4425, A1=>nx2256);
   ix2257 : xnor2 port map ( Y=>nx2256, A0=>nx4428, A1=>nx2254);
   ix4429 : aoi32 port map ( Y=>nx4428, A0=>nx5904, A1=>nx5900, A2=>nx2064, 
      B0=>nx1976, B1=>nx2066);
   ix2255 : xnor2 port map ( Y=>nx2254, A0=>nx4433, A1=>nx2252);
   ix2253 : xnor2 port map ( Y=>nx2252, A0=>nx4437, A1=>nx2250);
   ix4438 : aoi32 port map ( Y=>nx4437, A0=>nx5898, A1=>nx5908, A2=>nx2060, 
      B0=>nx1984, B1=>nx2062);
   ix2251 : xnor2 port map ( Y=>nx2250, A0=>nx4443, A1=>nx2248);
   ix2249 : xnor2 port map ( Y=>nx2248, A0=>nx4447, A1=>nx2246);
   ix4448 : aoi32 port map ( Y=>nx4447, A0=>nx5890, A1=>nx5916, A2=>nx2056, 
      B0=>nx1992, B1=>nx2058);
   ix2247 : xnor2 port map ( Y=>nx2246, A0=>nx4453, A1=>nx2244);
   ix2245 : xnor2 port map ( Y=>nx2244, A0=>nx4457, A1=>nx2242);
   ix4458 : aoi32 port map ( Y=>nx4457, A0=>nx5882, A1=>nx5924, A2=>nx2052, 
      B0=>nx2000, B1=>nx2054);
   ix2243 : xnor2 port map ( Y=>nx2242, A0=>nx4461, A1=>nx2240);
   ix2241 : xnor2 port map ( Y=>nx2240, A0=>nx4465, A1=>nx2238);
   ix4466 : aoi32 port map ( Y=>nx4465, A0=>nx5874, A1=>nx5932, A2=>nx2048, 
      B0=>nx2008, B1=>nx2050);
   ix2239 : xnor2 port map ( Y=>nx2238, A0=>nx4471, A1=>nx2236);
   ix2237 : xnor2 port map ( Y=>nx2236, A0=>nx4475, A1=>nx2234);
   ix4476 : aoi32 port map ( Y=>nx4475, A0=>nx5866, A1=>nx5940, A2=>nx2044, 
      B0=>nx2016, B1=>nx2046);
   ix2235 : xnor2 port map ( Y=>nx2234, A0=>nx4481, A1=>nx2232);
   ix2233 : xnor2 port map ( Y=>nx2232, A0=>nx2212, A1=>nx4493);
   ix2213 : oai32 port map ( Y=>nx2212, A0=>nx6020, A1=>nx6118, A2=>nx4335, 
      B0=>nx4487, B1=>nx4331);
   ix4494 : xnor2 port map ( Y=>nx4493, A0=>nx4495, A1=>nx4497);
   ix4498 : nand02 port map ( Y=>nx4497, A0=>nx5854, A1=>nx5964);
   MAC0_RegMultInB_reg_Y_15 : dffr port map ( Q=>OPEN, QB=>nx4503, D=>nx2222, 
      CLK=>clk, R=>nx5816);
   ix4508 : xnor2 port map ( Y=>nx4507, A0=>nx2783, A1=>nx4254);
   ix4255 : xnor2 port map ( Y=>nx4254, A0=>MAC0_adderB_15, A1=>
      RegOut_dup0_15);
   MAC0_RegMultOut_reg_Y_16 : dffr port map ( Q=>MAC0_adderB_16, QB=>OPEN, D
      =>nx3818, CLK=>clk, R=>nx5816);
   ix3819 : xnor2 port map ( Y=>nx3818, A0=>nx2300, A1=>nx4516);
   ix2301 : nor03 port map ( Y=>nx2300, A0=>nx4365, A1=>nx6132, A2=>nx6140);
   ix4518 : xnor2 port map ( Y=>nx4516, A0=>nx4519, A1=>nx4521);
   ix4522 : xnor2 port map ( Y=>nx4521, A0=>nx4523, A1=>nx4525);
   ix4524 : aoi32 port map ( Y=>nx4523, A0=>nx5960, A1=>nx5850, A2=>nx2280, 
      B0=>nx2108, B1=>nx2282);
   ix4526 : xnor2 port map ( Y=>nx4525, A0=>nx4527, A1=>nx4529);
   ix4530 : xnor2 port map ( Y=>nx4529, A0=>nx4531, A1=>nx4535);
   ix4532 : aoi32 port map ( Y=>nx4531, A0=>nx5952, A1=>nx5862, A2=>nx2276, 
      B0=>nx2116, B1=>nx2278);
   ix4536 : xnor2 port map ( Y=>nx4535, A0=>nx4537, A1=>nx4539);
   ix4540 : xnor2 port map ( Y=>nx4539, A0=>nx4541, A1=>nx4544);
   ix4542 : aoi32 port map ( Y=>nx4541, A0=>nx5944, A1=>nx5870, A2=>nx2272, 
      B0=>nx2124, B1=>nx2274);
   ix4545 : xnor2 port map ( Y=>nx4544, A0=>nx4547, A1=>nx4549);
   ix4550 : xnor2 port map ( Y=>nx4549, A0=>nx4551, A1=>nx4554);
   ix4552 : aoi32 port map ( Y=>nx4551, A0=>nx5936, A1=>nx5878, A2=>nx2268, 
      B0=>nx2132, B1=>nx2270);
   ix4556 : xnor2 port map ( Y=>nx4554, A0=>nx4557, A1=>nx4559);
   ix4560 : xnor2 port map ( Y=>nx4559, A0=>nx4561, A1=>nx4565);
   ix4562 : aoi32 port map ( Y=>nx4561, A0=>nx5928, A1=>nx5886, A2=>nx2264, 
      B0=>nx2140, B1=>nx2266);
   ix4566 : xnor2 port map ( Y=>nx4565, A0=>nx4567, A1=>nx4569);
   ix4570 : xnor2 port map ( Y=>nx4569, A0=>nx4571, A1=>nx4575);
   ix4572 : aoi32 port map ( Y=>nx4571, A0=>nx5920, A1=>nx5894, A2=>nx2260, 
      B0=>nx2148, B1=>nx2262);
   ix4576 : xnor2 port map ( Y=>nx4575, A0=>nx4577, A1=>nx4579);
   ix4580 : xnor2 port map ( Y=>nx4579, A0=>nx4581, A1=>nx4584);
   ix4582 : aoi32 port map ( Y=>nx4581, A0=>nx5912, A1=>nx5902, A2=>nx2256, 
      B0=>nx2156, B1=>nx2258);
   ix4585 : xnor2 port map ( Y=>nx4584, A0=>nx4587, A1=>nx4589);
   ix4590 : xnor2 port map ( Y=>nx4589, A0=>nx4591, A1=>nx4595);
   ix4592 : aoi32 port map ( Y=>nx4591, A0=>nx5906, A1=>nx5908, A2=>nx2252, 
      B0=>nx2164, B1=>nx2254);
   ix4596 : xnor2 port map ( Y=>nx4595, A0=>nx4597, A1=>nx4599);
   ix4600 : xnor2 port map ( Y=>nx4599, A0=>nx4601, A1=>nx4604);
   ix4602 : aoi32 port map ( Y=>nx4601, A0=>nx5898, A1=>nx5916, A2=>nx2248, 
      B0=>nx2172, B1=>nx2250);
   ix4605 : xnor2 port map ( Y=>nx4604, A0=>nx4607, A1=>nx4609);
   ix4610 : xnor2 port map ( Y=>nx4609, A0=>nx4611, A1=>nx4615);
   ix4612 : aoi32 port map ( Y=>nx4611, A0=>nx5890, A1=>nx5924, A2=>nx2244, 
      B0=>nx2180, B1=>nx2246);
   ix4616 : xnor2 port map ( Y=>nx4615, A0=>nx4617, A1=>nx4619);
   ix4620 : xnor2 port map ( Y=>nx4619, A0=>nx4621, A1=>nx4624);
   ix4622 : aoi32 port map ( Y=>nx4621, A0=>nx5882, A1=>nx5932, A2=>nx2240, 
      B0=>nx2188, B1=>nx2242);
   ix4625 : xnor2 port map ( Y=>nx4624, A0=>nx4627, A1=>nx4629);
   ix4630 : xnor2 port map ( Y=>nx4629, A0=>nx4631, A1=>nx4635);
   ix4632 : aoi32 port map ( Y=>nx4631, A0=>nx5874, A1=>nx5940, A2=>nx2236, 
      B0=>nx2196, B1=>nx2238);
   ix4636 : xnor2 port map ( Y=>nx4635, A0=>nx4637, A1=>nx4639);
   ix4640 : xnor2 port map ( Y=>nx4639, A0=>nx4641, A1=>nx4644);
   ix4642 : aoi32 port map ( Y=>nx4641, A0=>nx5866, A1=>nx5948, A2=>nx2232, 
      B0=>nx2204, B1=>nx2234);
   ix4645 : xnor2 port map ( Y=>nx4644, A0=>nx4647, A1=>nx4649);
   ix4650 : mux21 port map ( Y=>nx4649, A0=>nx4651, A1=>nx2414, S0=>nx2412);
   ix2415 : nor02 port map ( Y=>nx2414, A0=>nx6020, A1=>nx6136);
   ix2413 : oai32 port map ( Y=>nx2412, A0=>nx6020, A1=>nx6128, A2=>nx4497, 
      B0=>nx4656, B1=>nx4493);
   ix4666 : xnor2 port map ( Y=>nx4665, A0=>nx2775, A1=>nx4270);
   ix4271 : xnor2 port map ( Y=>nx4270, A0=>MAC0_adderB_16, A1=>
      RegOut_dup0_16);
   MAC0_RegMultOut_reg_Y_17 : dffr port map ( Q=>MAC0_adderB_17, QB=>OPEN, D
      =>nx3812, CLK=>clk, R=>nx5816);
   ix3813 : xor2 port map ( Y=>nx3812, A0=>nx2484, A1=>nx2644);
   ix2485 : oai32 port map ( Y=>nx2484, A0=>nx6132, A1=>nx6016, A2=>nx4521, 
      B0=>nx4674, B1=>nx4516);
   ix2645 : xnor2 port map ( Y=>nx2644, A0=>nx4677, A1=>nx2642);
   ix2643 : xnor2 port map ( Y=>nx2642, A0=>nx2492, A1=>nx4681);
   ix2493 : oai32 port map ( Y=>nx2492, A0=>nx6122, A1=>nx6030, A2=>nx4529, 
      B0=>nx4523, B1=>nx4525);
   ix4682 : xnor2 port map ( Y=>nx4681, A0=>nx4683, A1=>nx4685);
   ix4686 : xnor2 port map ( Y=>nx4685, A0=>nx2500, A1=>nx2636);
   ix2501 : oai32 port map ( Y=>nx2500, A0=>nx6114, A1=>nx6038, A2=>nx4539, 
      B0=>nx4531, B1=>nx4535);
   ix2637 : xnor2 port map ( Y=>nx2636, A0=>nx4689, A1=>nx2634);
   ix2635 : xnor2 port map ( Y=>nx2634, A0=>nx2508, A1=>nx4693);
   ix2509 : oai32 port map ( Y=>nx2508, A0=>nx6106, A1=>nx6046, A2=>nx4549, 
      B0=>nx4541, B1=>nx4544);
   ix4694 : xnor2 port map ( Y=>nx4693, A0=>nx4695, A1=>nx4697);
   ix4698 : xnor2 port map ( Y=>nx4697, A0=>nx2516, A1=>nx2628);
   ix2517 : oai32 port map ( Y=>nx2516, A0=>nx6098, A1=>nx6054, A2=>nx4559, 
      B0=>nx4551, B1=>nx4554);
   ix2629 : xnor2 port map ( Y=>nx2628, A0=>nx4701, A1=>nx2626);
   ix2627 : xnor2 port map ( Y=>nx2626, A0=>nx2524, A1=>nx4705);
   ix2525 : oai32 port map ( Y=>nx2524, A0=>nx6090, A1=>nx6062, A2=>nx4569, 
      B0=>nx4561, B1=>nx4565);
   ix4706 : xnor2 port map ( Y=>nx4705, A0=>nx4707, A1=>nx4709);
   ix4710 : xnor2 port map ( Y=>nx4709, A0=>nx2532, A1=>nx2620);
   ix2533 : oai32 port map ( Y=>nx2532, A0=>nx6082, A1=>nx6070, A2=>nx4579, 
      B0=>nx4571, B1=>nx4575);
   ix2621 : xnor2 port map ( Y=>nx2620, A0=>nx4713, A1=>nx2618);
   ix2619 : xnor2 port map ( Y=>nx2618, A0=>nx2540, A1=>nx4717);
   ix2541 : oai32 port map ( Y=>nx2540, A0=>nx6074, A1=>nx6078, A2=>nx4589, 
      B0=>nx4581, B1=>nx4584);
   ix4718 : xnor2 port map ( Y=>nx4717, A0=>nx4719, A1=>nx4721);
   ix4722 : xnor2 port map ( Y=>nx4721, A0=>nx2548, A1=>nx2612);
   ix2549 : oai32 port map ( Y=>nx2548, A0=>nx6066, A1=>nx6086, A2=>nx4599, 
      B0=>nx4591, B1=>nx4595);
   ix2613 : xnor2 port map ( Y=>nx2612, A0=>nx4725, A1=>nx2610);
   ix2611 : xnor2 port map ( Y=>nx2610, A0=>nx2556, A1=>nx4729);
   ix2557 : oai32 port map ( Y=>nx2556, A0=>nx6058, A1=>nx6094, A2=>nx4609, 
      B0=>nx4601, B1=>nx4604);
   ix4730 : xnor2 port map ( Y=>nx4729, A0=>nx4731, A1=>nx4733);
   ix4734 : xnor2 port map ( Y=>nx4733, A0=>nx2564, A1=>nx2604);
   ix2565 : oai32 port map ( Y=>nx2564, A0=>nx6050, A1=>nx6102, A2=>nx4619, 
      B0=>nx4611, B1=>nx4615);
   ix2605 : xnor2 port map ( Y=>nx2604, A0=>nx4737, A1=>nx2602);
   ix2603 : xnor2 port map ( Y=>nx2602, A0=>nx2572, A1=>nx4741);
   ix2573 : oai32 port map ( Y=>nx2572, A0=>nx6042, A1=>nx6110, A2=>nx4629, 
      B0=>nx4621, B1=>nx4624);
   ix4742 : xnor2 port map ( Y=>nx4741, A0=>nx4743, A1=>nx4745);
   ix4746 : xnor2 port map ( Y=>nx4745, A0=>nx2580, A1=>nx2596);
   ix2581 : oai32 port map ( Y=>nx2580, A0=>nx6034, A1=>nx6118, A2=>nx4639, 
      B0=>nx4631, B1=>nx4635);
   ix2597 : xnor2 port map ( Y=>nx2596, A0=>nx4749, A1=>nx2594);
   ix2595 : xnor2 port map ( Y=>nx2594, A0=>nx2588, A1=>nx4753);
   ix2589 : oai32 port map ( Y=>nx2588, A0=>nx6026, A1=>nx6128, A2=>nx4649, 
      B0=>nx4641, B1=>nx4644);
   ix4754 : xnor2 port map ( Y=>nx4753, A0=>nx4755, A1=>nx4757);
   ix4764 : xnor2 port map ( Y=>nx4763, A0=>nx2767, A1=>nx4286);
   ix4287 : xnor2 port map ( Y=>nx4286, A0=>MAC0_adderB_17, A1=>
      RegOut_dup0_17);
   MAC0_RegMultOut_reg_Y_18 : dffr port map ( Q=>MAC0_adderB_18, QB=>OPEN, D
      =>nx3806, CLK=>clk, R=>nx5816);
   ix3807 : xnor2 port map ( Y=>nx3806, A0=>nx4771, A1=>nx2804);
   ix4772 : aoi32 port map ( Y=>nx4771, A0=>nx5968, A1=>nx5862, A2=>nx2642, 
      B0=>nx2484, B1=>nx2644);
   ix2805 : xnor2 port map ( Y=>nx2804, A0=>nx4775, A1=>nx2802);
   ix2803 : xnor2 port map ( Y=>nx2802, A0=>nx2658, A1=>nx4781);
   ix2659 : oai32 port map ( Y=>nx2658, A0=>nx6122, A1=>nx6038, A2=>nx4685, 
      B0=>nx4779, B1=>nx4681);
   ix4780 : inv01 port map ( Y=>nx4779, A=>nx2492);
   ix4782 : xnor2 port map ( Y=>nx4781, A0=>nx4783, A1=>nx4785);
   ix4786 : xnor2 port map ( Y=>nx4785, A0=>nx4787, A1=>nx4789);
   ix4788 : aoi32 port map ( Y=>nx4787, A0=>nx5952, A1=>nx5878, A2=>nx2634, 
      B0=>nx2500, B1=>nx2636);
   ix4790 : xnor2 port map ( Y=>nx4789, A0=>nx4791, A1=>nx4793);
   ix4794 : xnor2 port map ( Y=>nx4793, A0=>nx2674, A1=>nx2792);
   ix2675 : oai32 port map ( Y=>nx2674, A0=>nx6106, A1=>nx6054, A2=>nx4697, 
      B0=>nx4797, B1=>nx4693);
   ix4798 : inv01 port map ( Y=>nx4797, A=>nx2508);
   ix2793 : xnor2 port map ( Y=>nx2792, A0=>nx4801, A1=>nx2790);
   ix2791 : xnor2 port map ( Y=>nx2790, A0=>nx4805, A1=>nx2788);
   ix4806 : aoi32 port map ( Y=>nx4805, A0=>nx5936, A1=>nx5894, A2=>nx2626, 
      B0=>nx2516, B1=>nx2628);
   ix2789 : xnor2 port map ( Y=>nx2788, A0=>nx4809, A1=>nx2786);
   ix2787 : xnor2 port map ( Y=>nx2786, A0=>nx2690, A1=>nx4817);
   ix2691 : oai32 port map ( Y=>nx2690, A0=>nx6090, A1=>nx6070, A2=>nx4709, 
      B0=>nx4815, B1=>nx4705);
   ix4816 : inv01 port map ( Y=>nx4815, A=>nx2524);
   ix4818 : xnor2 port map ( Y=>nx4817, A0=>nx4819, A1=>nx4821);
   ix4822 : xnor2 port map ( Y=>nx4821, A0=>nx4823, A1=>nx4825);
   ix4824 : aoi32 port map ( Y=>nx4823, A0=>nx5922, A1=>nx5910, A2=>nx2618, 
      B0=>nx2532, B1=>nx2620);
   ix4826 : xnor2 port map ( Y=>nx4825, A0=>nx4827, A1=>nx4829);
   ix4830 : xnor2 port map ( Y=>nx4829, A0=>nx2706, A1=>nx2776);
   ix2707 : oai32 port map ( Y=>nx2706, A0=>nx6074, A1=>nx6086, A2=>nx4721, 
      B0=>nx4833, B1=>nx4717);
   ix4834 : inv01 port map ( Y=>nx4833, A=>nx2540);
   ix2777 : xnor2 port map ( Y=>nx2776, A0=>nx4837, A1=>nx2774);
   ix2775 : xnor2 port map ( Y=>nx2774, A0=>nx4841, A1=>nx2772);
   ix4842 : aoi32 port map ( Y=>nx4841, A0=>nx5906, A1=>nx5924, A2=>nx2610, 
      B0=>nx2548, B1=>nx2612);
   ix2773 : xnor2 port map ( Y=>nx2772, A0=>nx4845, A1=>nx2770);
   ix2771 : xnor2 port map ( Y=>nx2770, A0=>nx2722, A1=>nx4853);
   ix2723 : oai32 port map ( Y=>nx2722, A0=>nx6058, A1=>nx6102, A2=>nx4733, 
      B0=>nx4851, B1=>nx4729);
   ix4852 : inv01 port map ( Y=>nx4851, A=>nx2556);
   ix4854 : xnor2 port map ( Y=>nx4853, A0=>nx4855, A1=>nx4857);
   ix4858 : xnor2 port map ( Y=>nx4857, A0=>nx4859, A1=>nx4861);
   ix4860 : aoi32 port map ( Y=>nx4859, A0=>nx5890, A1=>nx5940, A2=>nx2602, 
      B0=>nx2564, B1=>nx2604);
   ix4862 : xnor2 port map ( Y=>nx4861, A0=>nx4863, A1=>nx4865);
   ix4866 : xnor2 port map ( Y=>nx4865, A0=>nx2738, A1=>nx2760);
   ix2739 : oai32 port map ( Y=>nx2738, A0=>nx6042, A1=>nx6118, A2=>nx4745, 
      B0=>nx4869, B1=>nx4741);
   ix4870 : inv01 port map ( Y=>nx4869, A=>nx2572);
   ix2761 : xnor2 port map ( Y=>nx2760, A0=>nx4873, A1=>nx2758);
   ix2759 : xnor2 port map ( Y=>nx2758, A0=>nx4877, A1=>nx2756);
   ix4878 : aoi32 port map ( Y=>nx4877, A0=>nx5874, A1=>nx5956, A2=>nx2594, 
      B0=>nx2580, B1=>nx2596);
   ix2757 : xnor2 port map ( Y=>nx2756, A0=>nx4881, A1=>nx2754);
   ix2755 : oai32 port map ( Y=>nx2754, A0=>nx6026, A1=>nx6136, A2=>nx4757, 
      B0=>nx4884, B1=>nx4753);
   ix4885 : inv01 port map ( Y=>nx4884, A=>nx2588);
   ix4890 : xnor2 port map ( Y=>nx4889, A0=>nx2759, A1=>nx4302);
   ix4303 : xnor2 port map ( Y=>nx4302, A0=>MAC0_adderB_18, A1=>
      RegOut_dup0_18);
   MAC0_RegMultOut_reg_Y_19 : dffr port map ( Q=>MAC0_adderB_19, QB=>OPEN, D
      =>nx3800, CLK=>clk, R=>nx5818);
   ix3801 : xor2 port map ( Y=>nx3800, A0=>nx4896, A1=>nx4899);
   ix4897 : aoi32 port map ( Y=>nx4896, A0=>nx5968, A1=>nx5870, A2=>nx2802, 
      B0=>nx2650, B1=>nx2804);
   ix4900 : xnor2 port map ( Y=>nx4899, A0=>nx4901, A1=>nx4903);
   ix4904 : xnor2 port map ( Y=>nx4903, A0=>nx2818, A1=>nx2948);
   ix2819 : oai32 port map ( Y=>nx2818, A0=>nx6122, A1=>nx6046, A2=>nx4785, 
      B0=>nx4906, B1=>nx4781);
   ix2949 : xnor2 port map ( Y=>nx2948, A0=>nx4911, A1=>nx2946);
   ix2947 : xnor2 port map ( Y=>nx2946, A0=>nx2826, A1=>nx4915);
   ix2827 : oai32 port map ( Y=>nx2826, A0=>nx6114, A1=>nx6054, A2=>nx4793, 
      B0=>nx4787, B1=>nx4789);
   ix4916 : xnor2 port map ( Y=>nx4915, A0=>nx4917, A1=>nx4919);
   ix4920 : xnor2 port map ( Y=>nx4919, A0=>nx4921, A1=>nx4923);
   ix4922 : aoi32 port map ( Y=>nx4921, A0=>nx5944, A1=>nx5894, A2=>nx2790, 
      B0=>nx2674, B1=>nx2792);
   ix4924 : xnor2 port map ( Y=>nx4923, A0=>nx4925, A1=>nx4927);
   ix4928 : xnor2 port map ( Y=>nx4927, A0=>nx4929, A1=>nx4932);
   ix4930 : aoi32 port map ( Y=>nx4929, A0=>nx5936, A1=>nx5902, A2=>nx2786, 
      B0=>nx2682, B1=>nx2788);
   ix4933 : xnor2 port map ( Y=>nx4932, A0=>nx4934, A1=>nx4936);
   ix4937 : xnor2 port map ( Y=>nx4936, A0=>nx2850, A1=>nx2932);
   ix2851 : oai32 port map ( Y=>nx2850, A0=>nx6090, A1=>nx6078, A2=>nx4821, 
      B0=>nx4939, B1=>nx4817);
   ix2933 : xnor2 port map ( Y=>nx2932, A0=>nx4944, A1=>nx2930);
   ix2931 : xnor2 port map ( Y=>nx2930, A0=>nx2858, A1=>nx4948);
   ix2859 : oai32 port map ( Y=>nx2858, A0=>nx6082, A1=>nx6086, A2=>nx4829, 
      B0=>nx4823, B1=>nx4825);
   ix4949 : xnor2 port map ( Y=>nx4948, A0=>nx4950, A1=>nx4952);
   ix4953 : xnor2 port map ( Y=>nx4952, A0=>nx4954, A1=>nx4956);
   ix4955 : aoi32 port map ( Y=>nx4954, A0=>nx5914, A1=>nx5926, A2=>nx2774, 
      B0=>nx2706, B1=>nx2776);
   ix4957 : xnor2 port map ( Y=>nx4956, A0=>nx4958, A1=>nx4960);
   ix4961 : xnor2 port map ( Y=>nx4960, A0=>nx4962, A1=>nx4965);
   ix4963 : aoi32 port map ( Y=>nx4962, A0=>nx5906, A1=>nx5932, A2=>nx2770, 
      B0=>nx2714, B1=>nx2772);
   ix4966 : xnor2 port map ( Y=>nx4965, A0=>nx4967, A1=>nx4969);
   ix4970 : xnor2 port map ( Y=>nx4969, A0=>nx2882, A1=>nx2916);
   ix2883 : oai32 port map ( Y=>nx2882, A0=>nx6058, A1=>nx6110, A2=>nx4857, 
      B0=>nx4972, B1=>nx4853);
   ix2917 : xnor2 port map ( Y=>nx2916, A0=>nx4977, A1=>nx2914);
   ix2915 : xnor2 port map ( Y=>nx2914, A0=>nx2890, A1=>nx4981);
   ix2891 : oai32 port map ( Y=>nx2890, A0=>nx6050, A1=>nx6118, A2=>nx4865, 
      B0=>nx4859, B1=>nx4861);
   ix4982 : xnor2 port map ( Y=>nx4981, A0=>nx4983, A1=>nx4985);
   ix4986 : xnor2 port map ( Y=>nx4985, A0=>nx4987, A1=>nx4989);
   ix4988 : aoi32 port map ( Y=>nx4987, A0=>nx5882, A1=>nx5956, A2=>nx2758, 
      B0=>nx2738, B1=>nx2760);
   ix4990 : xnor2 port map ( Y=>nx4989, A0=>nx4991, A1=>nx4993);
   ix4994 : aoi32 port map ( Y=>nx4993, A0=>nx5874, A1=>nx5964, A2=>nx2754, 
      B0=>nx2746, B1=>nx2756);
   ix5000 : xnor2 port map ( Y=>nx4999, A0=>nx2751, A1=>nx4318);
   ix4319 : xnor2 port map ( Y=>nx4318, A0=>MAC0_adderB_19, A1=>
      RegOut_dup0_19);
   MAC0_RegMultOut_reg_Y_20 : dffr port map ( Q=>MAC0_adderB_20, QB=>OPEN, D
      =>nx3794, CLK=>clk, R=>nx5818);
   ix3795 : xnor2 port map ( Y=>nx3794, A0=>nx2958, A1=>nx5007);
   ix2959 : oai32 port map ( Y=>nx2958, A0=>nx6132, A1=>nx6046, A2=>nx4903, 
      B0=>nx4896, B1=>nx4899);
   ix5008 : xnor2 port map ( Y=>nx5007, A0=>nx5009, A1=>nx5011);
   ix5012 : xnor2 port map ( Y=>nx5011, A0=>nx5013, A1=>nx5015);
   ix5014 : aoi32 port map ( Y=>nx5013, A0=>nx5960, A1=>nx5886, A2=>nx2946, 
      B0=>nx2818, B1=>nx2948);
   ix5016 : xnor2 port map ( Y=>nx5015, A0=>nx5017, A1=>nx5019);
   ix5020 : xnor2 port map ( Y=>nx5019, A0=>nx2974, A1=>nx3080);
   ix2975 : oai32 port map ( Y=>nx2974, A0=>nx6114, A1=>nx6062, A2=>nx4919, 
      B0=>nx5022, B1=>nx4915);
   ix5023 : inv01 port map ( Y=>nx5022, A=>nx2826);
   ix3081 : xnor2 port map ( Y=>nx3080, A0=>nx5025, A1=>nx3078);
   ix3079 : xnor2 port map ( Y=>nx3078, A0=>nx2982, A1=>nx5029);
   ix2983 : oai32 port map ( Y=>nx2982, A0=>nx6106, A1=>nx6070, A2=>nx4927, 
      B0=>nx4921, B1=>nx4923);
   ix5030 : xnor2 port map ( Y=>nx5029, A0=>nx5031, A1=>nx5033);
   ix5034 : xnor2 port map ( Y=>nx5033, A0=>nx2990, A1=>nx3072);
   ix2991 : oai32 port map ( Y=>nx2990, A0=>nx6098, A1=>nx6078, A2=>nx4936, 
      B0=>nx4929, B1=>nx4932);
   ix3073 : xnor2 port map ( Y=>nx3072, A0=>nx5037, A1=>nx3070);
   ix3071 : xnor2 port map ( Y=>nx3070, A0=>nx5040, A1=>nx3068);
   ix5041 : aoi32 port map ( Y=>nx5040, A0=>nx5930, A1=>nx5918, A2=>nx2930, 
      B0=>nx2850, B1=>nx2932);
   ix3069 : xnor2 port map ( Y=>nx3068, A0=>nx5043, A1=>nx3066);
   ix3067 : xnor2 port map ( Y=>nx3066, A0=>nx3006, A1=>nx5049);
   ix3007 : oai32 port map ( Y=>nx3006, A0=>nx6082, A1=>nx6094, A2=>nx4952, 
      B0=>nx5047, B1=>nx4948);
   ix5048 : inv01 port map ( Y=>nx5047, A=>nx2858);
   ix5050 : xnor2 port map ( Y=>nx5049, A0=>nx5051, A1=>nx5053);
   ix5054 : xnor2 port map ( Y=>nx5053, A0=>nx3014, A1=>nx3060);
   ix3015 : oai32 port map ( Y=>nx3014, A0=>nx6074, A1=>nx6102, A2=>nx4960, 
      B0=>nx4954, B1=>nx4956);
   ix3061 : xnor2 port map ( Y=>nx3060, A0=>nx5057, A1=>nx3058);
   ix3059 : xnor2 port map ( Y=>nx3058, A0=>nx3022, A1=>nx5061);
   ix3023 : oai32 port map ( Y=>nx3022, A0=>nx6066, A1=>nx6110, A2=>nx4969, 
      B0=>nx4962, B1=>nx4965);
   ix5062 : xnor2 port map ( Y=>nx5061, A0=>nx5063, A1=>nx5065);
   ix5066 : xnor2 port map ( Y=>nx5065, A0=>nx5067, A1=>nx5069);
   ix5068 : aoi32 port map ( Y=>nx5067, A0=>nx5898, A1=>nx5948, A2=>nx2914, 
      B0=>nx2882, B1=>nx2916);
   ix5070 : xnor2 port map ( Y=>nx5069, A0=>nx5071, A1=>nx5073);
   ix5074 : xnor2 port map ( Y=>nx5073, A0=>nx3038, A1=>nx3048);
   ix3039 : oai32 port map ( Y=>nx3038, A0=>nx6050, A1=>nx6128, A2=>nx4985, 
      B0=>nx5076, B1=>nx4981);
   ix5077 : inv01 port map ( Y=>nx5076, A=>nx2890);
   ix3049 : xnor2 port map ( Y=>nx3048, A0=>nx5079, A1=>nx3046);
   ix3047 : oai32 port map ( Y=>nx3046, A0=>nx6042, A1=>nx6136, A2=>nx4993, 
      B0=>nx4987, B1=>nx4989);
   ix5086 : xnor2 port map ( Y=>nx5085, A0=>nx2743, A1=>nx4334);
   ix4335 : xnor2 port map ( Y=>nx4334, A0=>MAC0_adderB_20, A1=>
      RegOut_dup0_20);
   MAC0_RegMultOut_reg_Y_21 : dffr port map ( Q=>MAC0_adderB_21, QB=>OPEN, D
      =>nx3788, CLK=>clk, R=>nx5818);
   ix3789 : xor2 port map ( Y=>nx3788, A0=>nx3094, A1=>nx3212);
   ix3095 : oai32 port map ( Y=>nx3094, A0=>nx6132, A1=>nx6054, A2=>nx5011, 
      B0=>nx5093, B1=>nx5007);
   ix5094 : inv01 port map ( Y=>nx5093, A=>nx2958);
   ix3213 : xnor2 port map ( Y=>nx3212, A0=>nx5096, A1=>nx3210);
   ix3211 : xnor2 port map ( Y=>nx3210, A0=>nx3102, A1=>nx5100);
   ix3103 : oai32 port map ( Y=>nx3102, A0=>nx6122, A1=>nx6062, A2=>nx5019, 
      B0=>nx5013, B1=>nx5015);
   ix5101 : xnor2 port map ( Y=>nx5100, A0=>nx5102, A1=>nx5104);
   ix5105 : xnor2 port map ( Y=>nx5104, A0=>nx5106, A1=>nx5108);
   ix5107 : aoi32 port map ( Y=>nx5106, A0=>nx5952, A1=>nx5902, A2=>nx3078, 
      B0=>nx2974, B1=>nx3080);
   ix5109 : xnor2 port map ( Y=>nx5108, A0=>nx5110, A1=>nx5112);
   ix5113 : xnor2 port map ( Y=>nx5112, A0=>nx3118, A1=>nx3200);
   ix3119 : oai32 port map ( Y=>nx3118, A0=>nx6106, A1=>nx6078, A2=>nx5033, 
      B0=>nx5115, B1=>nx5029);
   ix5116 : inv01 port map ( Y=>nx5115, A=>nx2982);
   ix3201 : xnor2 port map ( Y=>nx3200, A0=>nx5118, A1=>nx3198);
   ix3199 : xnor2 port map ( Y=>nx3198, A0=>nx5121, A1=>nx3196);
   ix5122 : aoi32 port map ( Y=>nx5121, A0=>nx5938, A1=>nx5918, A2=>nx3070, 
      B0=>nx2990, B1=>nx3072);
   ix3197 : xnor2 port map ( Y=>nx3196, A0=>nx5124, A1=>nx3194);
   ix3195 : xnor2 port map ( Y=>nx3194, A0=>nx5127, A1=>nx3192);
   ix5128 : aoi32 port map ( Y=>nx5127, A0=>nx5930, A1=>nx5926, A2=>nx3066, 
      B0=>nx2998, B1=>nx3068);
   ix3193 : xnor2 port map ( Y=>nx3192, A0=>nx5131, A1=>nx3190);
   ix3191 : xnor2 port map ( Y=>nx3190, A0=>nx3142, A1=>nx5139);
   ix3143 : oai32 port map ( Y=>nx3142, A0=>nx6082, A1=>nx6102, A2=>nx5053, 
      B0=>nx5135, B1=>nx5049);
   ix5140 : xnor2 port map ( Y=>nx5139, A0=>nx5141, A1=>nx5143);
   ix5144 : xnor2 port map ( Y=>nx5143, A0=>nx5145, A1=>nx5147);
   ix5146 : aoi32 port map ( Y=>nx5145, A0=>nx5914, A1=>nx5940, A2=>nx3058, 
      B0=>nx3014, B1=>nx3060);
   ix5148 : xnor2 port map ( Y=>nx5147, A0=>nx5149, A1=>nx5151);
   ix5152 : xnor2 port map ( Y=>nx5151, A0=>nx3158, A1=>nx3180);
   ix3159 : oai32 port map ( Y=>nx3158, A0=>nx6066, A1=>nx6118, A2=>nx5065, 
      B0=>nx5154, B1=>nx5061);
   ix5155 : inv01 port map ( Y=>nx5154, A=>nx3022);
   ix3181 : xnor2 port map ( Y=>nx3180, A0=>nx5157, A1=>nx3178);
   ix3179 : xnor2 port map ( Y=>nx3178, A0=>nx3166, A1=>nx5161);
   ix3167 : oai32 port map ( Y=>nx3166, A0=>nx6058, A1=>nx6128, A2=>nx5073, 
      B0=>nx5067, B1=>nx5069);
   ix5162 : xnor2 port map ( Y=>nx5161, A0=>nx5163, A1=>nx5165);
   ix5166 : aoi32 port map ( Y=>nx5165, A0=>nx5890, A1=>nx5964, A2=>nx3046, 
      B0=>nx3038, B1=>nx3048);
   ix5171 : xnor2 port map ( Y=>nx5170, A0=>nx2735, A1=>nx4350);
   ix4351 : xnor2 port map ( Y=>nx4350, A0=>MAC0_adderB_21, A1=>
      RegOut_dup0_21);
   MAC0_RegMultOut_reg_Y_22 : dffr port map ( Q=>MAC0_adderB_22, QB=>OPEN, D
      =>nx3782, CLK=>clk, R=>nx5818);
   ix3783 : xnor2 port map ( Y=>nx3782, A0=>nx5177, A1=>nx3324);
   ix5178 : aoi32 port map ( Y=>nx5177, A0=>nx5968, A1=>nx5894, A2=>nx3210, 
      B0=>nx3094, B1=>nx3212);
   ix3325 : xnor2 port map ( Y=>nx3324, A0=>nx5180, A1=>nx3322);
   ix3323 : xnor2 port map ( Y=>nx3322, A0=>nx3226, A1=>nx5186);
   ix3227 : oai32 port map ( Y=>nx3226, A0=>nx6122, A1=>nx6070, A2=>nx5104, 
      B0=>nx5184, B1=>nx5100);
   ix5185 : inv01 port map ( Y=>nx5184, A=>nx3102);
   ix5187 : xnor2 port map ( Y=>nx5186, A0=>nx5188, A1=>nx5190);
   ix5191 : xnor2 port map ( Y=>nx5190, A0=>nx3234, A1=>nx3316);
   ix3235 : oai32 port map ( Y=>nx3234, A0=>nx6114, A1=>nx6078, A2=>nx5112, 
      B0=>nx5106, B1=>nx5108);
   ix3317 : xnor2 port map ( Y=>nx3316, A0=>nx5194, A1=>nx3314);
   ix3315 : xnor2 port map ( Y=>nx3314, A0=>nx5197, A1=>nx3312);
   ix5198 : aoi32 port map ( Y=>nx5197, A0=>nx5944, A1=>nx5918, A2=>nx3198, 
      B0=>nx3118, B1=>nx3200);
   ix3313 : xnor2 port map ( Y=>nx3312, A0=>nx5200, A1=>nx3310);
   ix3311 : xnor2 port map ( Y=>nx3310, A0=>nx5203, A1=>nx3308);
   ix5204 : aoi32 port map ( Y=>nx5203, A0=>nx5938, A1=>nx5926, A2=>nx3194, 
      B0=>nx3126, B1=>nx3196);
   ix3309 : xnor2 port map ( Y=>nx3308, A0=>nx5207, A1=>nx3306);
   ix3307 : xnor2 port map ( Y=>nx3306, A0=>nx5210, A1=>nx3304);
   ix5211 : aoi32 port map ( Y=>nx5210, A0=>nx5930, A1=>nx5934, A2=>nx3190, 
      B0=>nx3134, B1=>nx3192);
   ix3305 : xnor2 port map ( Y=>nx3304, A0=>nx5214, A1=>nx3302);
   ix3303 : xnor2 port map ( Y=>nx3302, A0=>nx3266, A1=>nx5222);
   ix3267 : oai32 port map ( Y=>nx3266, A0=>nx6082, A1=>nx6110, A2=>nx5143, 
      B0=>nx5218, B1=>nx5139);
   ix5223 : xnor2 port map ( Y=>nx5222, A0=>nx5224, A1=>nx5226);
   ix5227 : xnor2 port map ( Y=>nx5226, A0=>nx3274, A1=>nx3296);
   ix3275 : oai32 port map ( Y=>nx3274, A0=>nx6074, A1=>nx6118, A2=>nx5151, 
      B0=>nx5145, B1=>nx5147);
   ix3297 : xnor2 port map ( Y=>nx3296, A0=>nx5230, A1=>nx3294);
   ix3295 : xnor2 port map ( Y=>nx3294, A0=>nx5233, A1=>nx3292);
   ix5234 : aoi32 port map ( Y=>nx5233, A0=>nx5906, A1=>nx5956, A2=>nx3178, 
      B0=>nx3158, B1=>nx3180);
   ix3293 : xnor2 port map ( Y=>nx3292, A0=>nx5236, A1=>nx3290);
   ix3291 : oai32 port map ( Y=>nx3290, A0=>nx6058, A1=>nx6136, A2=>nx5165, 
      B0=>nx5239, B1=>nx5161);
   ix5240 : inv01 port map ( Y=>nx5239, A=>nx3166);
   ix5245 : xnor2 port map ( Y=>nx5244, A0=>nx2727, A1=>nx4366);
   ix4367 : xnor2 port map ( Y=>nx4366, A0=>MAC0_adderB_22, A1=>
      RegOut_dup0_22);
   MAC0_RegMultOut_reg_Y_23 : dffr port map ( Q=>MAC0_adderB_23, QB=>OPEN, D
      =>nx3776, CLK=>clk, R=>nx5818);
   ix3777 : xor2 port map ( Y=>nx3776, A0=>nx5251, A1=>nx5254);
   ix5252 : aoi32 port map ( Y=>nx5251, A0=>nx5968, A1=>nx5902, A2=>nx3322, 
      B0=>nx3218, B1=>nx3324);
   ix5255 : xnor2 port map ( Y=>nx5254, A0=>nx5256, A1=>nx5258);
   ix5259 : xnor2 port map ( Y=>nx5258, A0=>nx3338, A1=>nx3420);
   ix3339 : oai32 port map ( Y=>nx3338, A0=>nx6122, A1=>nx6078, A2=>nx5190, 
      B0=>nx5261, B1=>nx5186);
   ix3421 : xnor2 port map ( Y=>nx3420, A0=>nx5266, A1=>nx3418);
   ix3419 : xnor2 port map ( Y=>nx3418, A0=>nx5269, A1=>nx3416);
   ix5270 : aoi32 port map ( Y=>nx5269, A0=>nx5952, A1=>nx5918, A2=>nx3314, 
      B0=>nx3234, B1=>nx3316);
   ix3417 : xnor2 port map ( Y=>nx3416, A0=>nx5272, A1=>nx3414);
   ix3415 : xnor2 port map ( Y=>nx3414, A0=>nx5275, A1=>nx3412);
   ix5276 : aoi32 port map ( Y=>nx5275, A0=>nx5946, A1=>nx5926, A2=>nx3310, 
      B0=>nx3242, B1=>nx3312);
   ix3413 : xnor2 port map ( Y=>nx3412, A0=>nx5279, A1=>nx3410);
   ix3411 : xnor2 port map ( Y=>nx3410, A0=>nx5282, A1=>nx3408);
   ix5283 : aoi32 port map ( Y=>nx5282, A0=>nx5938, A1=>nx5934, A2=>nx3306, 
      B0=>nx3250, B1=>nx3308);
   ix3409 : xnor2 port map ( Y=>nx3408, A0=>nx5286, A1=>nx3406);
   ix3407 : xnor2 port map ( Y=>nx3406, A0=>nx5289, A1=>nx3404);
   ix5290 : aoi32 port map ( Y=>nx5289, A0=>nx5930, A1=>nx5942, A2=>nx3302, 
      B0=>nx3258, B1=>nx3304);
   ix3405 : xnor2 port map ( Y=>nx3404, A0=>nx5293, A1=>nx3402);
   ix3403 : xnor2 port map ( Y=>nx3402, A0=>nx3378, A1=>nx5301);
   ix3379 : oai32 port map ( Y=>nx3378, A0=>nx6082, A1=>nx6118, A2=>nx5226, 
      B0=>nx5297, B1=>nx5222);
   ix5302 : xnor2 port map ( Y=>nx5301, A0=>nx5303, A1=>nx5305);
   ix5306 : xnor2 port map ( Y=>nx5305, A0=>nx5307, A1=>nx5309);
   ix5308 : aoi32 port map ( Y=>nx5307, A0=>nx5914, A1=>nx5956, A2=>nx3294, 
      B0=>nx3274, B1=>nx3296);
   ix5310 : xnor2 port map ( Y=>nx5309, A0=>nx5311, A1=>nx5313);
   ix5314 : aoi32 port map ( Y=>nx5313, A0=>nx5906, A1=>nx5964, A2=>nx3290, 
      B0=>nx3282, B1=>nx3292);
   ix5320 : xnor2 port map ( Y=>nx5319, A0=>nx2719, A1=>nx4382);
   ix4383 : xnor2 port map ( Y=>nx4382, A0=>MAC0_adderB_23, A1=>
      RegOut_dup0_23);
   MAC0_RegMultOut_reg_Y_24 : dffr port map ( Q=>MAC0_adderB_24, QB=>OPEN, D
      =>nx3770, CLK=>clk, R=>nx5818);
   ix3771 : xnor2 port map ( Y=>nx3770, A0=>nx3430, A1=>nx5327);
   ix3431 : oai32 port map ( Y=>nx3430, A0=>nx6132, A1=>nx6078, A2=>nx5258, 
      B0=>nx5251, B1=>nx5254);
   ix5328 : xnor2 port map ( Y=>nx5327, A0=>nx5329, A1=>nx5331);
   ix5332 : xnor2 port map ( Y=>nx5331, A0=>nx5333, A1=>nx5335);
   ix5334 : aoi32 port map ( Y=>nx5333, A0=>nx5960, A1=>nx5918, A2=>nx3418, 
      B0=>nx3338, B1=>nx3420);
   ix5336 : xnor2 port map ( Y=>nx5335, A0=>nx5337, A1=>nx5339);
   ix5340 : xnor2 port map ( Y=>nx5339, A0=>nx5341, A1=>nx5344);
   ix5342 : aoi32 port map ( Y=>nx5341, A0=>nx5954, A1=>nx5926, A2=>nx3414, 
      B0=>nx3346, B1=>nx3416);
   ix5345 : xnor2 port map ( Y=>nx5344, A0=>nx5346, A1=>nx5348);
   ix5349 : xnor2 port map ( Y=>nx5348, A0=>nx5350, A1=>nx5353);
   ix5351 : aoi32 port map ( Y=>nx5350, A0=>nx5946, A1=>nx5934, A2=>nx3410, 
      B0=>nx3354, B1=>nx3412);
   ix5354 : xnor2 port map ( Y=>nx5353, A0=>nx5355, A1=>nx5357);
   ix5358 : xnor2 port map ( Y=>nx5357, A0=>nx5359, A1=>nx5362);
   ix5360 : aoi32 port map ( Y=>nx5359, A0=>nx5938, A1=>nx5942, A2=>nx3406, 
      B0=>nx3362, B1=>nx3408);
   ix5363 : xnor2 port map ( Y=>nx5362, A0=>nx5364, A1=>nx5366);
   ix5367 : xnor2 port map ( Y=>nx5366, A0=>nx5368, A1=>nx5371);
   ix5369 : aoi32 port map ( Y=>nx5368, A0=>nx5930, A1=>nx5948, A2=>nx3402, 
      B0=>nx3370, B1=>nx3404);
   ix5372 : xnor2 port map ( Y=>nx5371, A0=>nx5373, A1=>nx5375);
   ix5376 : xnor2 port map ( Y=>nx5375, A0=>nx3478, A1=>nx3488);
   ix3479 : oai32 port map ( Y=>nx3478, A0=>nx6082, A1=>nx6128, A2=>nx5305, 
      B0=>nx5378, B1=>nx5301);
   ix3489 : xnor2 port map ( Y=>nx3488, A0=>nx5383, A1=>nx3486);
   ix3487 : oai32 port map ( Y=>nx3486, A0=>nx6074, A1=>nx6136, A2=>nx5313, 
      B0=>nx5307, B1=>nx5309);
   ix5390 : xnor2 port map ( Y=>nx5389, A0=>nx2711, A1=>nx4398);
   ix4399 : xnor2 port map ( Y=>nx4398, A0=>MAC0_adderB_24, A1=>
      RegOut_dup0_24);
   MAC0_RegMultOut_reg_Y_25 : dffr port map ( Q=>MAC0_adderB_25, QB=>OPEN, D
      =>nx3764, CLK=>clk, R=>nx5818);
   ix3765 : xor2 port map ( Y=>nx3764, A0=>nx3518, A1=>nx3588);
   ix3519 : oai32 port map ( Y=>nx3518, A0=>nx6132, A1=>nx6086, A2=>nx5331, 
      B0=>nx5397, B1=>nx5327);
   ix5398 : inv01 port map ( Y=>nx5397, A=>nx3430);
   ix3589 : xnor2 port map ( Y=>nx3588, A0=>nx5400, A1=>nx3586);
   ix3587 : xnor2 port map ( Y=>nx3586, A0=>nx3526, A1=>nx5404);
   ix3527 : oai32 port map ( Y=>nx3526, A0=>nx6122, A1=>nx6094, A2=>nx5339, 
      B0=>nx5333, B1=>nx5335);
   ix5405 : xnor2 port map ( Y=>nx5404, A0=>nx5406, A1=>nx5408);
   ix5409 : xnor2 port map ( Y=>nx5408, A0=>nx3534, A1=>nx3580);
   ix3535 : oai32 port map ( Y=>nx3534, A0=>nx6114, A1=>nx6102, A2=>nx5348, 
      B0=>nx5341, B1=>nx5344);
   ix3581 : xnor2 port map ( Y=>nx3580, A0=>nx5412, A1=>nx3578);
   ix3579 : xnor2 port map ( Y=>nx3578, A0=>nx3542, A1=>nx5416);
   ix3543 : oai32 port map ( Y=>nx3542, A0=>nx6106, A1=>nx6110, A2=>nx5357, 
      B0=>nx5350, B1=>nx5353);
   ix5417 : xnor2 port map ( Y=>nx5416, A0=>nx5418, A1=>nx5420);
   ix5421 : xnor2 port map ( Y=>nx5420, A0=>nx3550, A1=>nx3572);
   ix3551 : oai32 port map ( Y=>nx3550, A0=>nx6098, A1=>nx6118, A2=>nx5366, 
      B0=>nx5359, B1=>nx5362);
   ix3573 : xnor2 port map ( Y=>nx3572, A0=>nx5424, A1=>nx3570);
   ix3571 : xnor2 port map ( Y=>nx3570, A0=>nx3558, A1=>nx5428);
   ix3559 : oai32 port map ( Y=>nx3558, A0=>nx6090, A1=>nx6128, A2=>nx5375, 
      B0=>nx5368, B1=>nx5371);
   ix5429 : xnor2 port map ( Y=>nx5428, A0=>nx5430, A1=>nx5432);
   ix5433 : aoi32 port map ( Y=>nx5432, A0=>nx5922, A1=>nx5966, A2=>nx3486, 
      B0=>nx3478, B1=>nx3488);
   ix5438 : xnor2 port map ( Y=>nx5437, A0=>nx2703, A1=>nx4414);
   ix4415 : xnor2 port map ( Y=>nx4414, A0=>MAC0_adderB_25, A1=>
      RegOut_dup0_25);
   MAC0_RegMultOut_reg_Y_26 : dffr port map ( Q=>MAC0_adderB_26, QB=>OPEN, D
      =>nx3758, CLK=>clk, R=>nx5820);
   ix3759 : xnor2 port map ( Y=>nx3758, A0=>nx5444, A1=>nx3652);
   ix5445 : aoi32 port map ( Y=>nx5444, A0=>nx5970, A1=>nx5926, A2=>nx3586, 
      B0=>nx3518, B1=>nx3588);
   ix3653 : xnor2 port map ( Y=>nx3652, A0=>nx5447, A1=>nx3650);
   ix3651 : xnor2 port map ( Y=>nx3650, A0=>nx3602, A1=>nx5453);
   ix3603 : oai32 port map ( Y=>nx3602, A0=>nx6122, A1=>nx6102, A2=>nx5408, 
      B0=>nx5451, B1=>nx5404);
   ix5452 : inv01 port map ( Y=>nx5451, A=>nx3526);
   ix5454 : xnor2 port map ( Y=>nx5453, A0=>nx5455, A1=>nx5457);
   ix5458 : xnor2 port map ( Y=>nx5457, A0=>nx5459, A1=>nx5461);
   ix5460 : aoi32 port map ( Y=>nx5459, A0=>nx5954, A1=>nx5942, A2=>nx3578, 
      B0=>nx3534, B1=>nx3580);
   ix5462 : xnor2 port map ( Y=>nx5461, A0=>nx5463, A1=>nx5465);
   ix5466 : xnor2 port map ( Y=>nx5465, A0=>nx3618, A1=>nx3640);
   ix3619 : oai32 port map ( Y=>nx3618, A0=>nx6106, A1=>nx6118, A2=>nx5420, 
      B0=>nx5468, B1=>nx5416);
   ix5469 : inv01 port map ( Y=>nx5468, A=>nx3542);
   ix3641 : xnor2 port map ( Y=>nx3640, A0=>nx5471, A1=>nx3638);
   ix3639 : xnor2 port map ( Y=>nx3638, A0=>nx5474, A1=>nx3636);
   ix5475 : aoi32 port map ( Y=>nx5474, A0=>nx5938, A1=>nx5958, A2=>nx3570, 
      B0=>nx3550, B1=>nx3572);
   ix3637 : xnor2 port map ( Y=>nx3636, A0=>nx5477, A1=>nx3634);
   ix3635 : oai32 port map ( Y=>nx3634, A0=>nx6090, A1=>nx6136, A2=>nx5432, 
      B0=>nx5480, B1=>nx5428);
   ix5481 : inv01 port map ( Y=>nx5480, A=>nx3558);
   ix5486 : xnor2 port map ( Y=>nx5485, A0=>nx2695, A1=>nx4430);
   ix4431 : xnor2 port map ( Y=>nx4430, A0=>MAC0_adderB_26, A1=>
      RegOut_dup0_26);
   MAC0_RegMultOut_reg_Y_27 : dffr port map ( Q=>MAC0_adderB_27, QB=>OPEN, D
      =>nx3752, CLK=>clk, R=>nx5820);
   ix3753 : xor2 port map ( Y=>nx3752, A0=>nx5492, A1=>nx5495);
   ix5493 : aoi32 port map ( Y=>nx5492, A0=>nx5970, A1=>nx5934, A2=>nx3650, 
      B0=>nx3594, B1=>nx3652);
   ix5496 : xnor2 port map ( Y=>nx5495, A0=>nx5497, A1=>nx5499);
   ix5500 : xnor2 port map ( Y=>nx5499, A0=>nx3666, A1=>nx3700);
   ix3667 : oai32 port map ( Y=>nx3666, A0=>nx6122, A1=>nx6110, A2=>nx5457, 
      B0=>nx5502, B1=>nx5453);
   ix3701 : xnor2 port map ( Y=>nx3700, A0=>nx5507, A1=>nx3698);
   ix3699 : xnor2 port map ( Y=>nx3698, A0=>nx3674, A1=>nx5511);
   ix3675 : oai32 port map ( Y=>nx3674, A0=>nx6114, A1=>nx6118, A2=>nx5465, 
      B0=>nx5459, B1=>nx5461);
   ix5512 : xnor2 port map ( Y=>nx5511, A0=>nx5513, A1=>nx5515);
   ix5516 : xnor2 port map ( Y=>nx5515, A0=>nx5517, A1=>nx5519);
   ix5518 : aoi32 port map ( Y=>nx5517, A0=>nx5946, A1=>nx5958, A2=>nx3638, 
      B0=>nx3618, B1=>nx3640);
   ix5520 : xnor2 port map ( Y=>nx5519, A0=>nx5521, A1=>nx5523);
   ix5524 : aoi32 port map ( Y=>nx5523, A0=>nx5938, A1=>nx5966, A2=>nx3634, 
      B0=>nx3626, B1=>nx3636);
   ix5530 : xnor2 port map ( Y=>nx5529, A0=>nx2687, A1=>nx4446);
   ix4447 : xnor2 port map ( Y=>nx4446, A0=>MAC0_adderB_27, A1=>
      RegOut_dup0_27);
   MAC0_RegMultOut_reg_Y_28 : dffr port map ( Q=>MAC0_adderB_28, QB=>OPEN, D
      =>nx3746, CLK=>clk, R=>nx5820);
   ix3747 : xnor2 port map ( Y=>nx3746, A0=>nx3710, A1=>nx5537);
   ix3711 : oai32 port map ( Y=>nx3710, A0=>nx6132, A1=>nx6110, A2=>nx5499, 
      B0=>nx5492, B1=>nx5495);
   ix5538 : xnor2 port map ( Y=>nx5537, A0=>nx5539, A1=>nx5541);
   ix5542 : xnor2 port map ( Y=>nx5541, A0=>nx5543, A1=>nx5545);
   ix5544 : aoi32 port map ( Y=>nx5543, A0=>nx5962, A1=>nx5950, A2=>nx3698, 
      B0=>nx3666, B1=>nx3700);
   ix5546 : xnor2 port map ( Y=>nx5545, A0=>nx5547, A1=>nx5549);
   ix5550 : xnor2 port map ( Y=>nx5549, A0=>nx3726, A1=>nx3736);
   ix3727 : oai32 port map ( Y=>nx3726, A0=>nx6114, A1=>nx6128, A2=>nx5515, 
      B0=>nx5552, B1=>nx5511);
   ix5553 : inv01 port map ( Y=>nx5552, A=>nx3674);
   ix3737 : xnor2 port map ( Y=>nx3736, A0=>nx5555, A1=>nx3734);
   ix3735 : oai32 port map ( Y=>nx3734, A0=>nx6106, A1=>nx6136, A2=>nx5523, 
      B0=>nx5517, B1=>nx5519);
   ix5562 : xnor2 port map ( Y=>nx5561, A0=>nx2679, A1=>nx4462);
   ix4463 : xnor2 port map ( Y=>nx4462, A0=>MAC0_adderB_28, A1=>
      RegOut_dup0_28);
   MAC0_RegMultOut_reg_Y_29 : dffr port map ( Q=>MAC0_adderB_29, QB=>OPEN, D
      =>nx4502, CLK=>clk, R=>nx5820);
   ix4503 : xor2 port map ( Y=>nx4502, A0=>nx4478, A1=>nx4500);
   ix4479 : oai32 port map ( Y=>nx4478, A0=>nx6132, A1=>nx6118, A2=>nx5541, 
      B0=>nx5569, B1=>nx5537);
   ix5570 : inv01 port map ( Y=>nx5569, A=>nx3710);
   ix4501 : xnor2 port map ( Y=>nx4500, A0=>nx5572, A1=>nx4498);
   ix4499 : xnor2 port map ( Y=>nx4498, A0=>nx4486, A1=>nx5576);
   ix4487 : oai32 port map ( Y=>nx4486, A0=>nx6122, A1=>nx6128, A2=>nx5549, 
      B0=>nx5543, B1=>nx5545);
   ix5577 : xnor2 port map ( Y=>nx5576, A0=>nx5578, A1=>nx5580);
   ix5581 : aoi32 port map ( Y=>nx5580, A0=>nx5954, A1=>nx5966, A2=>nx3734, 
      B0=>nx3726, B1=>nx3736);
   MISR0_reg_internal_reg_30 : dffr port map ( Q=>MISR_out_30, QB=>nx5584, D
      =>nx2309, CLK=>clk, R=>nx5820);
   MAC0_BigBoyReg_reg_Y_30 : dffr port map ( Q=>RegOut_dup0_30, QB=>OPEN, D
      =>nx1989, CLK=>clk, R=>nx5820);
   ix1990 : mux21 port map ( Y=>nx1989, A0=>RegOut_dup0_30, A1=>nx4548, S0=>
      WE);
   ix5593 : aoi22 port map ( Y=>nx5592, A0=>RegOut_dup0_29, A1=>nx4472, B0=>
      MAC0_adderB_29, B1=>nx5595);
   ix5596 : xnor2 port map ( Y=>nx5595, A0=>nx2671, A1=>nx4508);
   ix4509 : xnor2 port map ( Y=>nx4508, A0=>MAC0_adderB_29, A1=>
      RegOut_dup0_29);
   MAC0_RegMultOut_reg_Y_30 : dffr port map ( Q=>MAC0_adderB_30, QB=>OPEN, D
      =>nx4540, CLK=>clk, R=>nx5820);
   ix4541 : xnor2 port map ( Y=>nx4540, A0=>nx5602, A1=>nx4538);
   ix5603 : aoi32 port map ( Y=>nx5602, A0=>nx5970, A1=>nx5958, A2=>nx4498, 
      B0=>nx4478, B1=>nx4500);
   ix4539 : xnor2 port map ( Y=>nx4538, A0=>nx5605, A1=>nx4536);
   ix4537 : oai32 port map ( Y=>nx4536, A0=>nx6122, A1=>nx6136, A2=>nx5580, 
      B0=>nx5608, B1=>nx5576);
   ix5609 : inv01 port map ( Y=>nx5608, A=>nx4486);
   MISR0_reg_internal_reg_31 : dffr port map ( Q=>MISR_out_31, QB=>OPEN, D=>
      nx2299, CLK=>clk, R=>nx5820);
   MAC0_BigBoyReg_reg_Y_31 : dffr port map ( Q=>RegOut_dup0_31, QB=>OPEN, D
      =>nx1999, CLK=>clk, R=>nx5820);
   ix2000 : mux21 port map ( Y=>nx1999, A0=>RegOut_dup0_31, A1=>nx4574, S0=>
      WE);
   ix4575 : xnor2 port map ( Y=>nx4574, A0=>nx5620, A1=>nx5626);
   ix5621 : aoi22 port map ( Y=>nx5620, A0=>RegOut_dup0_30, A1=>nx4522, B0=>
      MAC0_adderB_30, B1=>nx5623);
   ix5624 : xnor2 port map ( Y=>nx5623, A0=>nx5592, A1=>nx4546);
   ix4547 : xnor2 port map ( Y=>nx4546, A0=>MAC0_adderB_30, A1=>
      RegOut_dup0_30);
   ix5627 : xor2 port map ( Y=>nx5626, A0=>MAC0_adderB_31, A1=>
      RegOut_dup0_31);
   MAC0_RegMultOut_reg_Y_31 : dffr port map ( Q=>MAC0_adderB_31, QB=>OPEN, D
      =>nx4566, CLK=>clk, R=>nx5820);
   MISR0_reg_internal_reg_0 : dffr port map ( Q=>MISR_out_0, QB=>nx5633, D=>
      nx2289, CLK=>clk, R=>nx5820);
   MISR0_reg_internal_reg_1 : dffr port map ( Q=>MISR_out_1, QB=>nx5638, D=>
      nx2279, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_2 : dffr port map ( Q=>MISR_out_2, QB=>nx5643, D=>
      nx2269, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_3 : dffs port map ( Q=>MISR_out_3, QB=>nx5648, D=>
      nx2259, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_4 : dffs port map ( Q=>MISR_out_4, QB=>nx5653, D=>
      nx2249, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_5 : dffs port map ( Q=>MISR_out_5, QB=>OPEN, D=>
      nx2239, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_6 : dffs port map ( Q=>MISR_out_6, QB=>OPEN, D=>
      nx2229, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_7 : dffr port map ( Q=>MISR_out_7, QB=>OPEN, D=>
      nx2219, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_8 : dffr port map ( Q=>MISR_out_8, QB=>OPEN, D=>
      nx2209, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_9 : dffs port map ( Q=>MISR_out_9, QB=>nx5678, D=>
      nx2199, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_10 : dffs port map ( Q=>MISR_out_10, QB=>nx5683, D
      =>nx2189, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_11 : dffr port map ( Q=>MISR_out_11, QB=>nx5688, D
      =>nx2179, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_12 : dffs port map ( Q=>MISR_out_12, QB=>nx5693, D
      =>nx2169, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_13 : dffr port map ( Q=>MISR_out_13, QB=>nx5698, D
      =>nx2159, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_14 : dffs port map ( Q=>MISR_out_14, QB=>nx5703, D
      =>nx2149, CLK=>clk, S=>nx5822);
   MISR0_reg_internal_reg_15 : dffr port map ( Q=>MISR_out_15, QB=>nx5708, D
      =>nx2139, CLK=>clk, R=>nx5822);
   MISR0_reg_internal_reg_16 : dffr port map ( Q=>MISR_out_16, QB=>nx5713, D
      =>nx2129, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_17 : dffr port map ( Q=>MISR_out_17, QB=>nx5718, D
      =>nx2119, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_18 : dffs port map ( Q=>MISR_out_18, QB=>nx5723, D
      =>nx2109, CLK=>clk, S=>nx5824);
   MISR0_reg_internal_reg_19 : dffr port map ( Q=>MISR_out_19, QB=>nx5728, D
      =>nx2099, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_20 : dffs port map ( Q=>MISR_out_20, QB=>nx5782, D
      =>nx2089, CLK=>clk, S=>nx5824);
   MISR0_reg_internal_reg_21 : dffs port map ( Q=>MISR_out_21, QB=>nx5738, D
      =>nx2079, CLK=>clk, S=>nx5824);
   MISR0_reg_internal_reg_22 : dffr port map ( Q=>MISR_out_22, QB=>nx5743, D
      =>nx2069, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_23 : dffr port map ( Q=>MISR_out_23, QB=>OPEN, D=>
      nx2059, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_24 : dffr port map ( Q=>MISR_out_24, QB=>nx5753, D
      =>nx2049, CLK=>clk, R=>nx5824);
   ix5759 : xnor2 port map ( Y=>nx5758, A0=>RegOut_dup0_24, A1=>MISR_out_25
   );
   MISR0_reg_internal_reg_25 : dffs port map ( Q=>MISR_out_25, QB=>OPEN, D=>
      nx2039, CLK=>clk, S=>nx5824);
   MISR0_reg_internal_reg_26 : dffr port map ( Q=>MISR_out_26, QB=>nx5780, D
      =>nx2029, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_27 : dffr port map ( Q=>MISR_out_27, QB=>OPEN, D=>
      nx2019, CLK=>clk, R=>nx5824);
   MISR0_reg_internal_reg_28 : dffs port map ( Q=>MISR_out_28, QB=>nx5773, D
      =>nx2009, CLK=>clk, S=>nx5824);
   MISR0_reg_internal_reg_29 : dffr port map ( Q=>MISR_out_29, QB=>nx5778, D
      =>nx2319, CLK=>clk, R=>nx5824);
   ix5789 : nand04 port map ( Y=>nx5788, A0=>nx4838, A1=>nx4848, A2=>nx4860, 
      A3=>nx4870);
   ix4549 : inv01 port map ( Y=>nx4548, A=>nx5623);
   ix4523 : inv01 port map ( Y=>nx4522, A=>nx5592);
   ix4511 : inv01 port map ( Y=>nx4510, A=>nx5595);
   ix4473 : inv01 port map ( Y=>nx4472, A=>nx2671);
   ix4465 : inv01 port map ( Y=>nx1041, A=>nx5561);
   ix4457 : inv01 port map ( Y=>nx4456, A=>nx2679);
   ix4449 : inv01 port map ( Y=>nx1039, A=>nx5529);
   ix4441 : inv01 port map ( Y=>nx4440, A=>nx2687);
   ix4433 : inv01 port map ( Y=>nx1037, A=>nx5485);
   ix4425 : inv01 port map ( Y=>nx4424, A=>nx2695);
   ix4417 : inv01 port map ( Y=>nx1035, A=>nx5437);
   ix4409 : inv01 port map ( Y=>nx4408, A=>nx2703);
   ix4401 : inv01 port map ( Y=>nx1033, A=>nx5389);
   ix4393 : inv01 port map ( Y=>nx4392, A=>nx2711);
   ix4385 : inv01 port map ( Y=>nx1031, A=>nx5319);
   ix4377 : inv01 port map ( Y=>nx4376, A=>nx2719);
   ix4369 : inv01 port map ( Y=>nx1029, A=>nx5244);
   ix4361 : inv01 port map ( Y=>nx4360, A=>nx2727);
   ix4353 : inv01 port map ( Y=>nx1027, A=>nx5170);
   ix4345 : inv01 port map ( Y=>nx4344, A=>nx2735);
   ix4337 : inv01 port map ( Y=>nx1025, A=>nx5085);
   ix4329 : inv01 port map ( Y=>nx4328, A=>nx2743);
   ix4321 : inv01 port map ( Y=>nx1023, A=>nx4999);
   ix4313 : inv01 port map ( Y=>nx4312, A=>nx2751);
   ix4305 : inv01 port map ( Y=>nx1021, A=>nx4889);
   ix4297 : inv01 port map ( Y=>nx4296, A=>nx2759);
   ix4289 : inv01 port map ( Y=>nx1019, A=>nx4763);
   ix4281 : inv01 port map ( Y=>nx4280, A=>nx2767);
   ix4273 : inv01 port map ( Y=>nx1017, A=>nx4665);
   ix4265 : inv01 port map ( Y=>nx4264, A=>nx2775);
   ix4257 : inv01 port map ( Y=>nx1015, A=>nx4507);
   ix4249 : inv01 port map ( Y=>nx4248, A=>nx2783);
   ix4241 : inv01 port map ( Y=>nx1013, A=>nx4347);
   ix4233 : inv01 port map ( Y=>nx4232, A=>nx2791);
   ix4225 : inv01 port map ( Y=>nx1011, A=>nx4201);
   ix4217 : inv01 port map ( Y=>nx4216, A=>nx2799);
   ix4209 : inv01 port map ( Y=>nx1009, A=>nx4061);
   ix4201 : inv01 port map ( Y=>nx4200, A=>nx2807);
   ix4193 : inv01 port map ( Y=>nx1007, A=>nx3939);
   ix4185 : inv01 port map ( Y=>nx4184, A=>nx2815);
   ix4177 : inv01 port map ( Y=>nx1005, A=>nx3823);
   ix4169 : inv01 port map ( Y=>nx4168, A=>nx2823);
   ix4161 : inv01 port map ( Y=>nx1003, A=>nx3725);
   ix4153 : inv01 port map ( Y=>nx4152, A=>nx2831);
   ix4145 : inv01 port map ( Y=>nx1001, A=>nx3615);
   ix4137 : inv01 port map ( Y=>nx4136, A=>nx2839);
   ix4129 : inv01 port map ( Y=>nx1000, A=>nx3515);
   ix4121 : inv01 port map ( Y=>nx4120, A=>nx2847);
   ix4113 : inv01 port map ( Y=>nx999, A=>nx3425);
   ix4105 : inv01 port map ( Y=>nx4104, A=>nx2855);
   ix4097 : inv01 port map ( Y=>nx998, A=>nx3347);
   ix4089 : inv01 port map ( Y=>nx4088, A=>nx2863);
   ix4081 : inv01 port map ( Y=>nx997, A=>nx3279);
   ix4073 : inv01 port map ( Y=>nx4072, A=>nx2871);
   ix4065 : inv01 port map ( Y=>nx995, A=>nx3225);
   ix4057 : inv01 port map ( Y=>nx4056, A=>nx2879);
   ix4049 : inv01 port map ( Y=>nx993, A=>nx3179);
   ix4041 : inv01 port map ( Y=>nx4040, A=>nx2887);
   ix4031 : inv01 port map ( Y=>nx991, A=>nx3143);
   ix3627 : inv01 port map ( Y=>nx3626, A=>nx5474);
   ix5503 : inv01 port map ( Y=>nx5502, A=>nx3602);
   ix3595 : inv01 port map ( Y=>nx3594, A=>nx5444);
   ix5379 : inv01 port map ( Y=>nx5378, A=>nx3378);
   ix3371 : inv01 port map ( Y=>nx3370, A=>nx5289);
   ix3363 : inv01 port map ( Y=>nx3362, A=>nx5282);
   ix3355 : inv01 port map ( Y=>nx3354, A=>nx5275);
   ix3347 : inv01 port map ( Y=>nx3346, A=>nx5269);
   ix3283 : inv01 port map ( Y=>nx3282, A=>nx5233);
   ix5298 : inv01 port map ( Y=>nx5297, A=>nx3266);
   ix3259 : inv01 port map ( Y=>nx3258, A=>nx5210);
   ix3251 : inv01 port map ( Y=>nx3250, A=>nx5203);
   ix3243 : inv01 port map ( Y=>nx3242, A=>nx5197);
   ix5262 : inv01 port map ( Y=>nx5261, A=>nx3226);
   ix3219 : inv01 port map ( Y=>nx3218, A=>nx5177);
   ix5219 : inv01 port map ( Y=>nx5218, A=>nx3142);
   ix3135 : inv01 port map ( Y=>nx3134, A=>nx5127);
   ix3127 : inv01 port map ( Y=>nx3126, A=>nx5121);
   ix5136 : inv01 port map ( Y=>nx5135, A=>nx3006);
   ix2999 : inv01 port map ( Y=>nx2998, A=>nx5040);
   ix2747 : inv01 port map ( Y=>nx2746, A=>nx4877);
   ix4973 : inv01 port map ( Y=>nx4972, A=>nx2722);
   ix2715 : inv01 port map ( Y=>nx2714, A=>nx4841);
   ix4940 : inv01 port map ( Y=>nx4939, A=>nx2690);
   ix2683 : inv01 port map ( Y=>nx2682, A=>nx4805);
   ix4907 : inv01 port map ( Y=>nx4906, A=>nx2658);
   ix2651 : inv01 port map ( Y=>nx2650, A=>nx4771);
   ix4675 : inv01 port map ( Y=>nx4674, A=>nx2300);
   ix4657 : inv01 port map ( Y=>nx4656, A=>nx2212);
   ix2205 : inv01 port map ( Y=>nx2204, A=>nx4475);
   ix2197 : inv01 port map ( Y=>nx2196, A=>nx4465);
   ix2189 : inv01 port map ( Y=>nx2188, A=>nx4457);
   ix2181 : inv01 port map ( Y=>nx2180, A=>nx4447);
   ix2173 : inv01 port map ( Y=>nx2172, A=>nx4437);
   ix2165 : inv01 port map ( Y=>nx2164, A=>nx4428);
   ix2157 : inv01 port map ( Y=>nx2156, A=>nx4419);
   ix2149 : inv01 port map ( Y=>nx2148, A=>nx4411);
   ix2141 : inv01 port map ( Y=>nx2140, A=>nx4401);
   ix2133 : inv01 port map ( Y=>nx2132, A=>nx4393);
   ix2125 : inv01 port map ( Y=>nx2124, A=>nx4383);
   ix2117 : inv01 port map ( Y=>nx2116, A=>nx4375);
   ix4488 : inv01 port map ( Y=>nx4487, A=>nx2024);
   ix2017 : inv01 port map ( Y=>nx2016, A=>nx4315);
   ix2009 : inv01 port map ( Y=>nx2008, A=>nx4305);
   ix2001 : inv01 port map ( Y=>nx2000, A=>nx4297);
   ix1993 : inv01 port map ( Y=>nx1992, A=>nx4287);
   ix1985 : inv01 port map ( Y=>nx1984, A=>nx4277);
   ix1977 : inv01 port map ( Y=>nx1976, A=>nx4268);
   ix1969 : inv01 port map ( Y=>nx1968, A=>nx4259);
   ix1961 : inv01 port map ( Y=>nx1960, A=>nx4251);
   ix1953 : inv01 port map ( Y=>nx1952, A=>nx4241);
   ix1945 : inv01 port map ( Y=>nx1944, A=>nx4233);
   ix1937 : inv01 port map ( Y=>nx1936, A=>nx4225);
   ix4326 : inv01 port map ( Y=>nx4325, A=>nx1848);
   ix1841 : inv01 port map ( Y=>nx1840, A=>nx4169);
   ix1833 : inv01 port map ( Y=>nx1832, A=>nx4159);
   ix1825 : inv01 port map ( Y=>nx1824, A=>nx4149);
   ix1817 : inv01 port map ( Y=>nx1816, A=>nx4140);
   ix1809 : inv01 port map ( Y=>nx1808, A=>nx4131);
   ix1801 : inv01 port map ( Y=>nx1800, A=>nx4123);
   ix1793 : inv01 port map ( Y=>nx1792, A=>nx4113);
   ix1785 : inv01 port map ( Y=>nx1784, A=>nx4105);
   ix1777 : inv01 port map ( Y=>nx1776, A=>nx4095);
   ix1769 : inv01 port map ( Y=>nx1768, A=>nx4089);
   ix4180 : inv01 port map ( Y=>nx4179, A=>nx1684);
   ix1677 : inv01 port map ( Y=>nx1676, A=>nx4031);
   ix1669 : inv01 port map ( Y=>nx1668, A=>nx4023);
   ix1661 : inv01 port map ( Y=>nx1660, A=>nx4015);
   ix1653 : inv01 port map ( Y=>nx1652, A=>nx4007);
   ix1645 : inv01 port map ( Y=>nx1644, A=>nx3999);
   ix1637 : inv01 port map ( Y=>nx1636, A=>nx3990);
   ix1629 : inv01 port map ( Y=>nx1628, A=>nx3981);
   ix1621 : inv01 port map ( Y=>nx1620, A=>nx3973);
   ix1613 : inv01 port map ( Y=>nx1612, A=>nx3965);
   ix4044 : inv01 port map ( Y=>nx4043, A=>nx1532);
   ix1525 : inv01 port map ( Y=>nx1524, A=>nx3909);
   ix1517 : inv01 port map ( Y=>nx1516, A=>nx3899);
   ix1509 : inv01 port map ( Y=>nx1508, A=>nx3891);
   ix1501 : inv01 port map ( Y=>nx1500, A=>nx3882);
   ix1493 : inv01 port map ( Y=>nx1492, A=>nx3873);
   ix1485 : inv01 port map ( Y=>nx1484, A=>nx3865);
   ix1477 : inv01 port map ( Y=>nx1476, A=>nx3857);
   ix1469 : inv01 port map ( Y=>nx1468, A=>nx3849);
   ix3920 : inv01 port map ( Y=>nx3919, A=>nx1392);
   ix1385 : inv01 port map ( Y=>nx1384, A=>nx3798);
   ix1377 : inv01 port map ( Y=>nx1376, A=>nx3791);
   ix1369 : inv01 port map ( Y=>nx1368, A=>nx3783);
   ix1361 : inv01 port map ( Y=>nx1360, A=>nx3774);
   ix1353 : inv01 port map ( Y=>nx1352, A=>nx3767);
   ix1345 : inv01 port map ( Y=>nx1344, A=>nx3759);
   ix1337 : inv01 port map ( Y=>nx1336, A=>nx3753);
   ix3808 : inv01 port map ( Y=>nx3807, A=>nx1264);
   ix1257 : inv01 port map ( Y=>nx1256, A=>nx3691);
   ix1249 : inv01 port map ( Y=>nx1248, A=>nx3681);
   ix1241 : inv01 port map ( Y=>nx1240, A=>nx3671);
   ix1233 : inv01 port map ( Y=>nx1232, A=>nx3661);
   ix1225 : inv01 port map ( Y=>nx1224, A=>nx3651);
   ix1217 : inv01 port map ( Y=>nx1216, A=>nx3643);
   ix3704 : inv01 port map ( Y=>nx3703, A=>nx1148);
   ix1141 : inv01 port map ( Y=>nx1140, A=>nx3581);
   ix1133 : inv01 port map ( Y=>nx1132, A=>nx3571);
   ix1125 : inv01 port map ( Y=>nx1124, A=>nx3561);
   ix1117 : inv01 port map ( Y=>nx1116, A=>nx3551);
   ix1109 : inv01 port map ( Y=>nx1108, A=>nx3543);
   ix3594 : inv01 port map ( Y=>nx3593, A=>nx1044);
   ix1037 : inv01 port map ( Y=>nx1036, A=>nx3481);
   ix1029 : inv01 port map ( Y=>nx1028, A=>nx3471);
   ix1021 : inv01 port map ( Y=>nx1020, A=>nx3461);
   ix1013 : inv01 port map ( Y=>nx1012, A=>nx3453);
   ix3494 : inv01 port map ( Y=>nx3493, A=>nx952);
   ix945 : inv01 port map ( Y=>nx944, A=>nx3391);
   ix937 : inv01 port map ( Y=>nx936, A=>nx3381);
   ix929 : inv01 port map ( Y=>nx928, A=>nx3373);
   ix3404 : inv01 port map ( Y=>nx3403, A=>nx872);
   ix865 : inv01 port map ( Y=>nx864, A=>nx3313);
   ix857 : inv01 port map ( Y=>nx856, A=>nx3305);
   ix3326 : inv01 port map ( Y=>nx3325, A=>nx804);
   ix797 : inv01 port map ( Y=>nx796, A=>nx3251);
   ix3262 : inv01 port map ( Y=>nx3261, A=>nx748);
   ix705 : inv01 port map ( Y=>nx704, A=>nx3207);
   ix5799 : inv02 port map ( Y=>nx5800, A=>reset);
   ix5801 : inv02 port map ( Y=>nx5802, A=>reset);
   ix5803 : inv02 port map ( Y=>nx5804, A=>reset);
   ix5805 : inv02 port map ( Y=>nx5806, A=>reset);
   ix5807 : inv02 port map ( Y=>nx5808, A=>reset);
   ix5809 : inv02 port map ( Y=>nx5810, A=>reset);
   ix5811 : inv02 port map ( Y=>nx5812, A=>reset);
   ix5813 : inv02 port map ( Y=>nx5814, A=>reset);
   ix5815 : inv02 port map ( Y=>nx5816, A=>reset);
   ix5817 : inv02 port map ( Y=>nx5818, A=>reset);
   ix5819 : inv02 port map ( Y=>nx5820, A=>reset);
   ix5821 : inv02 port map ( Y=>nx5822, A=>reset);
   ix5823 : inv02 port map ( Y=>nx5824, A=>reset);
   ix5843 : inv01 port map ( Y=>nx5844, A=>nx3135);
   ix5847 : inv01 port map ( Y=>nx5848, A=>nx3131);
   ix5849 : inv01 port map ( Y=>nx5850, A=>nx6016);
   ix5851 : buf02 port map ( Y=>nx5852, A=>MAC0_MultA_0);
   ix5853 : buf02 port map ( Y=>nx5854, A=>MAC0_MultA_0);
   ix5855 : inv01 port map ( Y=>nx5856, A=>nx6140);
   ix5859 : inv01 port map ( Y=>nx5860, A=>nx3173);
   ix5861 : inv01 port map ( Y=>nx5862, A=>nx6030);
   ix5863 : inv01 port map ( Y=>nx5864, A=>nx3159);
   ix5865 : inv01 port map ( Y=>nx5866, A=>nx6026);
   ix5867 : inv01 port map ( Y=>nx5868, A=>nx3219);
   ix5869 : inv01 port map ( Y=>nx5870, A=>nx6038);
   ix5871 : inv01 port map ( Y=>nx5872, A=>nx3195);
   ix5873 : inv01 port map ( Y=>nx5874, A=>nx6034);
   ix5875 : inv01 port map ( Y=>nx5876, A=>nx3273);
   ix5877 : inv01 port map ( Y=>nx5878, A=>nx6046);
   ix5879 : inv01 port map ( Y=>nx5880, A=>nx3241);
   ix5881 : inv01 port map ( Y=>nx5882, A=>nx6042);
   ix5883 : inv01 port map ( Y=>nx5884, A=>nx3341);
   ix5885 : inv01 port map ( Y=>nx5886, A=>nx6054);
   ix5887 : inv01 port map ( Y=>nx5888, A=>nx3295);
   ix5889 : inv01 port map ( Y=>nx5890, A=>nx6050);
   ix5891 : inv01 port map ( Y=>nx5892, A=>nx3419);
   ix5893 : inv01 port map ( Y=>nx5894, A=>nx6062);
   ix5895 : inv01 port map ( Y=>nx5896, A=>nx3363);
   ix5897 : inv01 port map ( Y=>nx5898, A=>nx6058);
   ix5899 : inv01 port map ( Y=>nx5900, A=>nx3509);
   ix5901 : inv01 port map ( Y=>nx5902, A=>nx6070);
   ix5903 : inv01 port map ( Y=>nx5904, A=>nx3441);
   ix5905 : inv01 port map ( Y=>nx5906, A=>nx6066);
   ix5907 : inv01 port map ( Y=>nx5908, A=>nx3609);
   ix5909 : inv01 port map ( Y=>nx5910, A=>nx6078);
   ix5911 : inv01 port map ( Y=>nx5912, A=>nx3531);
   ix5913 : inv01 port map ( Y=>nx5914, A=>nx6074);
   ix5915 : inv01 port map ( Y=>nx5916, A=>nx3719);
   ix5917 : inv01 port map ( Y=>nx5918, A=>nx6086);
   ix5919 : inv01 port map ( Y=>nx5920, A=>nx3631);
   ix5921 : inv01 port map ( Y=>nx5922, A=>nx6082);
   ix5923 : inv01 port map ( Y=>nx5924, A=>nx3819);
   ix5925 : inv01 port map ( Y=>nx5926, A=>nx6094);
   ix5927 : inv01 port map ( Y=>nx5928, A=>nx3741);
   ix5929 : inv01 port map ( Y=>nx5930, A=>nx6090);
   ix5931 : inv01 port map ( Y=>nx5932, A=>nx3933);
   ix5933 : inv01 port map ( Y=>nx5934, A=>nx6102);
   ix5935 : inv01 port map ( Y=>nx5936, A=>nx3837);
   ix5937 : inv01 port map ( Y=>nx5938, A=>nx6098);
   ix5939 : inv01 port map ( Y=>nx5940, A=>nx4057);
   ix5941 : inv01 port map ( Y=>nx5942, A=>nx6110);
   ix5943 : inv01 port map ( Y=>nx5944, A=>nx3953);
   ix5945 : inv01 port map ( Y=>nx5946, A=>nx6106);
   ix5947 : inv01 port map ( Y=>nx5948, A=>nx4195);
   ix5949 : inv01 port map ( Y=>nx5950, A=>nx6118);
   ix5951 : inv01 port map ( Y=>nx5952, A=>nx4076);
   ix5953 : inv01 port map ( Y=>nx5954, A=>nx6114);
   ix5955 : inv01 port map ( Y=>nx5956, A=>nx4341);
   ix5957 : inv01 port map ( Y=>nx5958, A=>nx6128);
   ix5959 : inv01 port map ( Y=>nx5960, A=>nx4215);
   ix5961 : inv01 port map ( Y=>nx5962, A=>nx6122);
   ix5963 : inv01 port map ( Y=>nx5964, A=>nx4503);
   ix5965 : inv01 port map ( Y=>nx5966, A=>nx6136);
   ix5967 : inv01 port map ( Y=>nx5968, A=>nx4363);
   ix5969 : inv01 port map ( Y=>nx5970, A=>nx6132);
   ix5971 : inv02 port map ( Y=>nx5972, A=>MAC0_MultB_0);
   ix5973 : inv02 port map ( Y=>nx5974, A=>MAC0_MultB_0);
   ix505 : or04 port map ( Y=>nx504, A0=>CounterOut_0, A1=>CounterOut_1, A2
      =>CounterOut_2, A3=>nx5980);
   ix5979 : inv01 port map ( Y=>nx5980, A=>CounterOut_3);
   ix1050 : xor2 port map ( Y=>nx1049, A0=>nx2339, A1=>nx5998);
   ix25 : or02 port map ( Y=>nx987, A0=>nx2339, A1=>nx2349);
   ix1070 : mux21 port map ( Y=>nx1069, A0=>nx30, A1=>CounterOut_2, S0=>
      nx5998);
   ix31 : xor2 port map ( Y=>nx30, A0=>nx987, A1=>nx2361);
   ix1080 : mux21 port map ( Y=>nx1079, A0=>nx44, A1=>CounterOut_3, S0=>
      nx5998);
   ix39 : or03 port map ( Y=>nx985, A0=>nx2339, A1=>nx2349, A2=>nx2361);
   ix497 : or04 port map ( Y=>nx496, A0=>CounterOut_4, A1=>nx2397, A2=>
      nx2407, A3=>nx2415);
   ix1090 : mux21 port map ( Y=>nx1089, A0=>nx58, A1=>CounterOut_4, S0=>
      nx5998);
   ix53 : or04 port map ( Y=>nx983, A0=>nx2339, A1=>nx2349, A2=>nx2361, A3=>
      nx5980);
   ix2390 : nor02ii port map ( Y=>nx2389, A0=>nx983, A1=>CounterOut_4);
   ix1100 : mux21 port map ( Y=>nx1099, A0=>nx72, A1=>CounterOut_5, S0=>
      nx5998);
   ix73 : xor2 port map ( Y=>nx72, A0=>nx2389, A1=>CounterOut_5);
   ix1110 : mux21 port map ( Y=>nx1109, A0=>nx86, A1=>CounterOut_6, S0=>
      nx5998);
   ix87 : xor2 port map ( Y=>nx86, A0=>nx979, A1=>nx2407);
   ix1120 : mux21 port map ( Y=>nx1119, A0=>nx100, A1=>CounterOut_7, S0=>
      nx5998);
   ix101 : xor2 port map ( Y=>nx100, A0=>nx2413, A1=>CounterOut_7);
   ix2414 : nor02ii port map ( Y=>nx2413, A0=>nx979, A1=>CounterOut_6);
   ix1130 : mux21 port map ( Y=>nx1129, A0=>nx114, A1=>CounterOut_8, S0=>
      nx5998);
   ix115 : xor2 port map ( Y=>nx114, A0=>nx975, A1=>nx2427);
   ix1140 : mux21 port map ( Y=>nx1139, A0=>nx128, A1=>CounterOut_9, S0=>
      nx5998);
   ix129 : xor2 port map ( Y=>nx128, A0=>nx2433, A1=>CounterOut_9);
   ix2434 : nor02ii port map ( Y=>nx2433, A0=>nx975, A1=>CounterOut_8);
   ix2438 : and02 port map ( Y=>nx2437, A0=>nx2447, A1=>nx2455);
   ix1150 : mux21 port map ( Y=>nx1149, A0=>nx142, A1=>CounterOut_10, S0=>
      nx5998);
   ix143 : xor2 port map ( Y=>nx142, A0=>nx971, A1=>nx2447);
   ix1160 : mux21 port map ( Y=>nx1159, A0=>nx156, A1=>CounterOut_11, S0=>
      nx5998);
   ix157 : xor2 port map ( Y=>nx156, A0=>nx2453, A1=>CounterOut_11);
   ix2454 : nor02ii port map ( Y=>nx2453, A0=>nx971, A1=>CounterOut_10);
   ix2458 : and04 port map ( Y=>nx2457, A0=>nx2467, A1=>nx2475, A2=>nx2485, 
      A3=>nx2493);
   ix1170 : mux21 port map ( Y=>nx1169, A0=>nx170, A1=>CounterOut_12, S0=>
      nx5998);
   ix171 : xor2 port map ( Y=>nx170, A0=>nx967, A1=>nx2467);
   ix1180 : mux21 port map ( Y=>nx1179, A0=>nx184, A1=>CounterOut_13, S0=>
      nx5998);
   ix185 : xor2 port map ( Y=>nx184, A0=>nx2473, A1=>CounterOut_13);
   ix2474 : nor02ii port map ( Y=>nx2473, A0=>nx967, A1=>CounterOut_12);
   ix1190 : mux21 port map ( Y=>nx1189, A0=>nx198, A1=>CounterOut_14, S0=>
      nx6000);
   ix199 : xor2 port map ( Y=>nx198, A0=>nx965, A1=>nx2485);
   ix1200 : mux21 port map ( Y=>nx1199, A0=>nx212, A1=>CounterOut_15, S0=>
      nx6000);
   ix213 : xor2 port map ( Y=>nx212, A0=>nx2491, A1=>CounterOut_15);
   ix2492 : nor02ii port map ( Y=>nx2491, A0=>nx965, A1=>CounterOut_14);
   ix2498 : and04 port map ( Y=>nx2497, A0=>nx2507, A1=>nx2515, A2=>nx2525, 
      A3=>nx2533);
   ix1210 : mux21 port map ( Y=>nx1209, A0=>nx226, A1=>CounterOut_16, S0=>
      nx6000);
   ix227 : xor2 port map ( Y=>nx226, A0=>nx963, A1=>nx2507);
   ix1220 : mux21 port map ( Y=>nx1219, A0=>nx240, A1=>CounterOut_17, S0=>
      nx6000);
   ix241 : xor2 port map ( Y=>nx240, A0=>nx2513, A1=>CounterOut_17);
   ix2514 : nor02ii port map ( Y=>nx2513, A0=>nx963, A1=>CounterOut_16);
   ix1230 : mux21 port map ( Y=>nx1229, A0=>nx254, A1=>CounterOut_18, S0=>
      nx6000);
   ix255 : xor2 port map ( Y=>nx254, A0=>nx959, A1=>nx2525);
   ix1240 : mux21 port map ( Y=>nx1239, A0=>nx268, A1=>CounterOut_19, S0=>
      nx6000);
   ix269 : xor2 port map ( Y=>nx268, A0=>nx2531, A1=>CounterOut_19);
   ix2532 : nor02ii port map ( Y=>nx2531, A0=>nx959, A1=>CounterOut_18);
   ix2536 : and04 port map ( Y=>nx2535, A0=>nx2545, A1=>nx2553, A2=>nx2563, 
      A3=>nx2571);
   ix1250 : mux21 port map ( Y=>nx1249, A0=>nx282, A1=>CounterOut_20, S0=>
      nx6000);
   ix283 : xor2 port map ( Y=>nx282, A0=>nx955, A1=>nx2545);
   ix1260 : mux21 port map ( Y=>nx1259, A0=>nx296, A1=>CounterOut_21, S0=>
      nx6000);
   ix297 : xor2 port map ( Y=>nx296, A0=>nx2551, A1=>CounterOut_21);
   ix2552 : nor02ii port map ( Y=>nx2551, A0=>nx955, A1=>CounterOut_20);
   ix1270 : mux21 port map ( Y=>nx1269, A0=>nx310, A1=>CounterOut_22, S0=>
      nx6000);
   ix311 : xor2 port map ( Y=>nx310, A0=>nx951, A1=>nx2563);
   ix1280 : mux21 port map ( Y=>nx1279, A0=>nx324, A1=>CounterOut_23, S0=>
      nx6000);
   ix325 : xor2 port map ( Y=>nx324, A0=>nx2569, A1=>CounterOut_23);
   ix2570 : nor02ii port map ( Y=>nx2569, A0=>nx951, A1=>CounterOut_22);
   ix2574 : and04 port map ( Y=>nx2573, A0=>nx2583, A1=>nx2591, A2=>nx2601, 
      A3=>nx2609);
   ix1290 : mux21 port map ( Y=>nx1289, A0=>nx338, A1=>CounterOut_24, S0=>
      nx6000);
   ix339 : xor2 port map ( Y=>nx338, A0=>nx947, A1=>nx2583);
   ix1300 : mux21 port map ( Y=>nx1299, A0=>nx352, A1=>CounterOut_25, S0=>
      nx6000);
   ix353 : xor2 port map ( Y=>nx352, A0=>nx2589, A1=>CounterOut_25);
   ix2590 : nor02ii port map ( Y=>nx2589, A0=>nx947, A1=>CounterOut_24);
   ix1310 : mux21 port map ( Y=>nx1309, A0=>nx366, A1=>CounterOut_26, S0=>
      nx6000);
   ix367 : xor2 port map ( Y=>nx366, A0=>nx943, A1=>nx2601);
   ix1320 : mux21 port map ( Y=>nx1319, A0=>nx380, A1=>CounterOut_27, S0=>
      nx6000);
   ix381 : xor2 port map ( Y=>nx380, A0=>nx2607, A1=>CounterOut_27);
   ix2608 : nor02ii port map ( Y=>nx2607, A0=>nx943, A1=>CounterOut_26);
   ix2612 : and04 port map ( Y=>nx2611, A0=>nx2621, A1=>nx2629, A2=>nx2639, 
      A3=>nx5982);
   ix5981 : inv01 port map ( Y=>nx5982, A=>CounterOut_31);
   ix1330 : mux21 port map ( Y=>nx1329, A0=>nx394, A1=>CounterOut_28, S0=>
      nx6000);
   ix395 : xor2 port map ( Y=>nx394, A0=>nx939, A1=>nx2621);
   ix1340 : mux21 port map ( Y=>nx1339, A0=>nx408, A1=>CounterOut_29, S0=>
      nx6002);
   ix409 : xor2 port map ( Y=>nx408, A0=>nx2627, A1=>CounterOut_29);
   ix2628 : nor02ii port map ( Y=>nx2627, A0=>nx939, A1=>CounterOut_28);
   ix1350 : mux21 port map ( Y=>nx1349, A0=>nx422, A1=>CounterOut_30, S0=>
      nx6002);
   ix423 : xor2 port map ( Y=>nx422, A0=>nx935, A1=>nx2639);
   ix1360 : mux21 port map ( Y=>nx1359, A0=>nx432, A1=>CounterOut_31, S0=>
      nx6002);
   ix2646 : nor02ii port map ( Y=>nx2645, A0=>nx935, A1=>CounterOut_30);
   ix4785 : and03 port map ( Y=>nx4784, A0=>nx5778, A1=>MISR_out_31, A2=>
      nx5584);
   ix2320 : mux21 port map ( Y=>nx2319, A0=>nx4772, A1=>MISR_out_29, S0=>
      nx6002);
   ix4773 : xor2 port map ( Y=>nx4772, A0=>RegOut_dup0_29, A1=>MISR_out_30);
   ix687 : mux21 port map ( Y=>nx686, A0=>LFSROUT_16, A1=>A(0), S0=>nx6002);
   ix1370 : mux21 port map ( Y=>nx1369, A0=>LFSROUT_17, A1=>LFSROUT_16, S0=>
      nx6002);
   ix1680 : mux21 port map ( Y=>nx1679, A0=>LFSROUT_18, A1=>LFSROUT_17, S0=>
      nx6002);
   ix1670 : mux21 port map ( Y=>nx1669, A0=>LFSROUT_19, A1=>LFSROUT_18, S0=>
      nx6002);
   ix1660 : mux21 port map ( Y=>nx1659, A0=>nx644, A1=>LFSROUT_19, S0=>
      nx6002);
   ix645 : xor2 port map ( Y=>nx644, A0=>LFSROUT_20, A1=>LFSROUT_0);
   ix1650 : mux21 port map ( Y=>nx1649, A0=>LFSROUT_21, A1=>LFSROUT_20, S0=>
      nx6002);
   ix1640 : mux21 port map ( Y=>nx1639, A0=>LFSROUT_22, A1=>LFSROUT_21, S0=>
      nx6002);
   ix1630 : mux21 port map ( Y=>nx1629, A0=>LFSROUT_23, A1=>LFSROUT_22, S0=>
      nx6002);
   ix1620 : mux21 port map ( Y=>nx1619, A0=>LFSROUT_24, A1=>LFSROUT_23, S0=>
      nx6002);
   ix1610 : mux21 port map ( Y=>nx1609, A0=>nx622, A1=>LFSROUT_24, S0=>
      nx6002);
   ix623 : xor2 port map ( Y=>nx622, A0=>LFSROUT_25, A1=>LFSROUT_0);
   ix1600 : mux21 port map ( Y=>nx1599, A0=>nx616, A1=>LFSROUT_25, S0=>
      nx6002);
   ix617 : xor2 port map ( Y=>nx616, A0=>LFSROUT_26, A1=>LFSROUT_0);
   ix1590 : mux21 port map ( Y=>nx1589, A0=>LFSROUT_27, A1=>LFSROUT_26, S0=>
      nx6004);
   ix1580 : mux21 port map ( Y=>nx1579, A0=>LFSROUT_28, A1=>LFSROUT_27, S0=>
      nx6004);
   ix1570 : mux21 port map ( Y=>nx1569, A0=>LFSROUT_29, A1=>LFSROUT_28, S0=>
      nx6004);
   ix1560 : mux21 port map ( Y=>nx1559, A0=>LFSROUT_30, A1=>LFSROUT_29, S0=>
      nx6004);
   ix1550 : mux21 port map ( Y=>nx1549, A0=>LFSROUT_31, A1=>LFSROUT_30, S0=>
      nx6004);
   ix1540 : mux21 port map ( Y=>nx1539, A0=>LFSROUT_0, A1=>LFSROUT_31, S0=>
      nx6004);
   ix1530 : mux21 port map ( Y=>nx1529, A0=>LFSROUT_1, A1=>LFSROUT_0, S0=>
      nx6004);
   ix1520 : mux21 port map ( Y=>nx1519, A0=>LFSROUT_2, A1=>LFSROUT_1, S0=>
      nx6004);
   ix1510 : mux21 port map ( Y=>nx1509, A0=>LFSROUT_3, A1=>LFSROUT_2, S0=>
      nx6004);
   ix1500 : mux21 port map ( Y=>nx1499, A0=>LFSROUT_4, A1=>LFSROUT_3, S0=>
      nx6004);
   ix1490 : mux21 port map ( Y=>nx1489, A0=>LFSROUT_5, A1=>LFSROUT_4, S0=>
      nx6004);
   ix1480 : mux21 port map ( Y=>nx1479, A0=>LFSROUT_6, A1=>LFSROUT_5, S0=>
      nx6004);
   ix1470 : mux21 port map ( Y=>nx1469, A0=>LFSROUT_7, A1=>LFSROUT_6, S0=>
      nx6004);
   ix1460 : mux21 port map ( Y=>nx1459, A0=>LFSROUT_8, A1=>LFSROUT_7, S0=>
      nx6004);
   ix1450 : mux21 port map ( Y=>nx1449, A0=>LFSROUT_9, A1=>LFSROUT_8, S0=>
      nx6004);
   ix1440 : mux21 port map ( Y=>nx1439, A0=>LFSROUT_10, A1=>LFSROUT_9, S0=>
      nx6006);
   ix1430 : mux21 port map ( Y=>nx1429, A0=>LFSROUT_11, A1=>LFSROUT_10, S0=>
      nx6006);
   ix1420 : mux21 port map ( Y=>nx1419, A0=>LFSROUT_12, A1=>LFSROUT_11, S0=>
      nx6006);
   ix1410 : mux21 port map ( Y=>nx1409, A0=>LFSROUT_13, A1=>LFSROUT_12, S0=>
      nx6006);
   ix1400 : mux21 port map ( Y=>nx1399, A0=>LFSROUT_14, A1=>LFSROUT_13, S0=>
      nx6006);
   ix1390 : mux21 port map ( Y=>nx1389, A0=>LFSROUT_15, A1=>LFSROUT_14, S0=>
      nx6006);
   ix1380 : mux21 port map ( Y=>nx1379, A0=>LFSROUT_16, A1=>LFSROUT_15, S0=>
      nx6006);
   ix699 : mux21 port map ( Y=>nx698, A0=>LFSROUT_0, A1=>B(0), S0=>nx6006);
   ix673 : mux21 port map ( Y=>nx672, A0=>LFSROUT_1, A1=>B(1), S0=>nx6006);
   ix661 : mux21 port map ( Y=>nx660, A0=>LFSROUT_17, A1=>A(1), S0=>nx6006);
   ix3138 : or04 port map ( Y=>nx3137, A0=>nx6020, A1=>nx6016, A2=>nx5984, 
      A3=>nx6140);
   ix5983 : inv01 port map ( Y=>nx5984, A=>nx5852);
   ix3154 : or02 port map ( Y=>nx3153, A0=>nx6026, A1=>nx6140);
   ix733 : mux21 port map ( Y=>nx732, A0=>LFSROUT_18, A1=>A(2), S0=>nx6006);
   ix3166 : or02 port map ( Y=>nx3165, A0=>nx6022, A1=>nx6016);
   ix715 : mux21 port map ( Y=>nx714, A0=>LFSROUT_2, A1=>B(2), S0=>nx6006);
   ix3190 : or02 port map ( Y=>nx3189, A0=>nx6034, A1=>nx6140);
   ix781 : mux21 port map ( Y=>nx780, A0=>LFSROUT_19, A1=>A(3), S0=>nx6006);
   ix3202 : or02 port map ( Y=>nx3201, A0=>nx6026, A1=>nx6016);
   ix3212 : or02 port map ( Y=>nx3211, A0=>nx6022, A1=>nx6030);
   ix759 : mux21 port map ( Y=>nx758, A0=>LFSROUT_3, A1=>B(3), S0=>nx6006);
   ix3236 : or02 port map ( Y=>nx3235, A0=>nx6042, A1=>nx6140);
   ix841 : mux21 port map ( Y=>nx840, A0=>LFSROUT_20, A1=>A(4), S0=>nx6006);
   ix3248 : or02 port map ( Y=>nx3247, A0=>nx6034, A1=>nx6016);
   ix3256 : or02 port map ( Y=>nx3255, A0=>nx6026, A1=>nx6030);
   ix3266 : or02 port map ( Y=>nx3265, A0=>nx6022, A1=>nx6038);
   ix815 : mux21 port map ( Y=>nx814, A0=>LFSROUT_4, A1=>B(4), S0=>nx6008);
   ix3290 : or02 port map ( Y=>nx3289, A0=>nx6050, A1=>nx6140);
   ix913 : mux21 port map ( Y=>nx912, A0=>LFSROUT_21, A1=>A(5), S0=>nx6008);
   ix3302 : or02 port map ( Y=>nx3301, A0=>nx6042, A1=>nx6016);
   ix3310 : or02 port map ( Y=>nx3309, A0=>nx6034, A1=>nx6030);
   ix3320 : or02 port map ( Y=>nx3319, A0=>nx6026, A1=>nx6038);
   ix3334 : or02 port map ( Y=>nx3333, A0=>nx6022, A1=>nx6046);
   ix883 : mux21 port map ( Y=>nx882, A0=>LFSROUT_5, A1=>B(5), S0=>nx6008);
   ix3358 : or02 port map ( Y=>nx3357, A0=>nx6058, A1=>nx6140);
   ix997 : mux21 port map ( Y=>nx996, A0=>LFSROUT_22, A1=>A(6), S0=>nx6008);
   ix3933 : nor02ii port map ( Y=>nx3932, A0=>nx6058, A1=>MAC0_MultB_0);
   ix3370 : or02 port map ( Y=>nx3369, A0=>nx6050, A1=>nx6016);
   ix3378 : or02 port map ( Y=>nx3377, A0=>nx6042, A1=>nx6030);
   ix3388 : or02 port map ( Y=>nx3387, A0=>nx6034, A1=>nx6038);
   ix3398 : or02 port map ( Y=>nx3397, A0=>nx6026, A1=>nx6046);
   ix3412 : or02 port map ( Y=>nx3411, A0=>nx6022, A1=>nx6054);
   ix963 : mux21 port map ( Y=>nx962, A0=>LFSROUT_6, A1=>B(6), S0=>nx6008);
   ix3436 : or02 port map ( Y=>nx3435, A0=>nx6066, A1=>nx6140);
   ix1093 : mux21 port map ( Y=>nx1092, A0=>LFSROUT_23, A1=>A(7), S0=>nx6008
   );
   ix3921 : nor02ii port map ( Y=>nx3920, A0=>nx6066, A1=>MAC0_MultB_0);
   ix3450 : or02 port map ( Y=>nx3449, A0=>nx6058, A1=>nx6016);
   ix3458 : or02 port map ( Y=>nx3457, A0=>nx6050, A1=>nx6030);
   ix3468 : or02 port map ( Y=>nx3467, A0=>nx6042, A1=>nx6038);
   ix3478 : or02 port map ( Y=>nx3477, A0=>nx6034, A1=>nx6046);
   ix3488 : or02 port map ( Y=>nx3487, A0=>nx6026, A1=>nx6054);
   ix3502 : or02 port map ( Y=>nx3501, A0=>nx6022, A1=>nx6062);
   ix1055 : mux21 port map ( Y=>nx1054, A0=>LFSROUT_7, A1=>B(7), S0=>nx6008
   );
   ix3526 : or02 port map ( Y=>nx3525, A0=>nx6074, A1=>nx6140);
   ix1201 : mux21 port map ( Y=>nx1200, A0=>LFSROUT_24, A1=>A(8), S0=>nx6008
   );
   ix3909 : nor02ii port map ( Y=>nx3908, A0=>nx6074, A1=>MAC0_MultB_0);
   ix3540 : or02 port map ( Y=>nx3539, A0=>nx6066, A1=>nx6016);
   ix3548 : or02 port map ( Y=>nx3547, A0=>nx6058, A1=>nx6030);
   ix3558 : or02 port map ( Y=>nx3557, A0=>nx6050, A1=>nx6038);
   ix3568 : or02 port map ( Y=>nx3567, A0=>nx6042, A1=>nx6046);
   ix3578 : or02 port map ( Y=>nx3577, A0=>nx6034, A1=>nx6054);
   ix3588 : or02 port map ( Y=>nx3587, A0=>nx6026, A1=>nx6062);
   ix3602 : or02 port map ( Y=>nx3601, A0=>nx6022, A1=>nx6070);
   ix1159 : mux21 port map ( Y=>nx1158, A0=>LFSROUT_8, A1=>B(8), S0=>nx6008
   );
   ix3626 : or02 port map ( Y=>nx3625, A0=>nx6082, A1=>nx6140);
   ix1321 : mux21 port map ( Y=>nx1320, A0=>LFSROUT_25, A1=>A(9), S0=>nx6008
   );
   ix3897 : nor02ii port map ( Y=>nx3896, A0=>nx6082, A1=>MAC0_MultB_0);
   ix3640 : or02 port map ( Y=>nx3639, A0=>nx6074, A1=>nx6016);
   ix3648 : or02 port map ( Y=>nx3647, A0=>nx6066, A1=>nx6030);
   ix3658 : or02 port map ( Y=>nx3657, A0=>nx6058, A1=>nx6038);
   ix3668 : or02 port map ( Y=>nx3667, A0=>nx6050, A1=>nx6046);
   ix3678 : or02 port map ( Y=>nx3677, A0=>nx6042, A1=>nx6054);
   ix3688 : or02 port map ( Y=>nx3687, A0=>nx6034, A1=>nx6062);
   ix3698 : or02 port map ( Y=>nx3697, A0=>nx6026, A1=>nx6070);
   ix3712 : or02 port map ( Y=>nx3711, A0=>nx6022, A1=>nx6078);
   ix1275 : mux21 port map ( Y=>nx1274, A0=>LFSROUT_9, A1=>B(9), S0=>nx6008
   );
   ix3736 : or02 port map ( Y=>nx3735, A0=>nx6090, A1=>nx5974);
   ix1453 : mux21 port map ( Y=>nx1452, A0=>LFSROUT_26, A1=>A(10), S0=>
      nx6008);
   ix3885 : nor02ii port map ( Y=>nx3884, A0=>nx6090, A1=>MAC0_MultB_0);
   ix3750 : or02 port map ( Y=>nx3749, A0=>nx6082, A1=>nx6016);
   ix3757 : or02 port map ( Y=>nx3756, A0=>nx6074, A1=>nx6030);
   ix3764 : or02 port map ( Y=>nx3763, A0=>nx6066, A1=>nx6038);
   ix3772 : or02 port map ( Y=>nx3771, A0=>nx6058, A1=>nx6046);
   ix3780 : or02 port map ( Y=>nx3779, A0=>nx6050, A1=>nx6054);
   ix3788 : or02 port map ( Y=>nx3787, A0=>nx6042, A1=>nx6062);
   ix3796 : or02 port map ( Y=>nx3795, A0=>nx6034, A1=>nx6070);
   ix3804 : or02 port map ( Y=>nx3803, A0=>nx6026, A1=>nx6078);
   ix3814 : or02 port map ( Y=>nx3813, A0=>nx6022, A1=>nx6086);
   ix1403 : mux21 port map ( Y=>nx1402, A0=>LFSROUT_10, A1=>B(10), S0=>
      nx6008);
   ix3834 : or02 port map ( Y=>nx3833, A0=>nx6098, A1=>nx5974);
   ix1597 : mux21 port map ( Y=>nx1596, A0=>LFSROUT_27, A1=>A(11), S0=>
      nx6008);
   ix3873 : nor02ii port map ( Y=>nx3872, A0=>nx6098, A1=>MAC0_MultB_0);
   ix3846 : or02 port map ( Y=>nx3845, A0=>nx6090, A1=>nx6016);
   ix3854 : or02 port map ( Y=>nx3853, A0=>nx6082, A1=>nx6030);
   ix3862 : or02 port map ( Y=>nx3861, A0=>nx6074, A1=>nx6038);
   ix3871 : or02 port map ( Y=>nx3870, A0=>nx6066, A1=>nx6046);
   ix3880 : or02 port map ( Y=>nx3879, A0=>nx6058, A1=>nx6054);
   ix3888 : or02 port map ( Y=>nx3887, A0=>nx6050, A1=>nx6062);
   ix3896 : or02 port map ( Y=>nx3895, A0=>nx6042, A1=>nx6070);
   ix3906 : or02 port map ( Y=>nx3905, A0=>nx6034, A1=>nx6078);
   ix3916 : or02 port map ( Y=>nx3915, A0=>nx6026, A1=>nx6086);
   ix3928 : or02 port map ( Y=>nx3927, A0=>nx6022, A1=>nx6094);
   ix1543 : mux21 port map ( Y=>nx1542, A0=>LFSROUT_11, A1=>B(11), S0=>
      nx6008);
   ix3948 : or02 port map ( Y=>nx3947, A0=>nx6106, A1=>nx5974);
   ix1753 : mux21 port map ( Y=>nx1752, A0=>LFSROUT_28, A1=>A(12), S0=>
      nx6010);
   ix3861 : nor02ii port map ( Y=>nx3860, A0=>nx6106, A1=>MAC0_MultB_0);
   ix3962 : or02 port map ( Y=>nx3961, A0=>nx6098, A1=>nx6016);
   ix3970 : or02 port map ( Y=>nx3969, A0=>nx6090, A1=>nx6030);
   ix3979 : or02 port map ( Y=>nx3978, A0=>nx6082, A1=>nx6038);
   ix3988 : or02 port map ( Y=>nx3987, A0=>nx6074, A1=>nx6046);
   ix3996 : or02 port map ( Y=>nx3995, A0=>nx6066, A1=>nx6054);
   ix4005 : or02 port map ( Y=>nx4004, A0=>nx6058, A1=>nx6062);
   ix4012 : or02 port map ( Y=>nx4011, A0=>nx6050, A1=>nx6070);
   ix4020 : or02 port map ( Y=>nx4019, A0=>nx6042, A1=>nx6078);
   ix4028 : or02 port map ( Y=>nx4027, A0=>nx6034, A1=>nx6086);
   ix4038 : or02 port map ( Y=>nx4037, A0=>nx6026, A1=>nx6094);
   ix4050 : or02 port map ( Y=>nx4049, A0=>nx6022, A1=>nx6102);
   ix1695 : mux21 port map ( Y=>nx1694, A0=>LFSROUT_12, A1=>B(12), S0=>
      nx6010);
   ix4072 : or02 port map ( Y=>nx4071, A0=>nx6114, A1=>nx5974);
   ix1921 : mux21 port map ( Y=>nx1920, A0=>LFSROUT_29, A1=>A(13), S0=>
      nx6010);
   ix3849 : nor02ii port map ( Y=>nx3848, A0=>nx6114, A1=>MAC0_MultB_0);
   ix4086 : or02 port map ( Y=>nx4085, A0=>nx6106, A1=>nx6016);
   ix4093 : or02 port map ( Y=>nx4092, A0=>nx6098, A1=>nx6030);
   ix4102 : or02 port map ( Y=>nx4101, A0=>nx6090, A1=>nx6038);
   ix4110 : or02 port map ( Y=>nx4109, A0=>nx6082, A1=>nx6046);
   ix4120 : or02 port map ( Y=>nx4119, A0=>nx6074, A1=>nx6054);
   ix4128 : or02 port map ( Y=>nx4127, A0=>nx6066, A1=>nx6062);
   ix4138 : or02 port map ( Y=>nx4137, A0=>nx6060, A1=>nx6070);
   ix4146 : or02 port map ( Y=>nx4145, A0=>nx6050, A1=>nx6078);
   ix4156 : or02 port map ( Y=>nx4155, A0=>nx6042, A1=>nx6086);
   ix4166 : or02 port map ( Y=>nx4165, A0=>nx6034, A1=>nx6094);
   ix4174 : or02 port map ( Y=>nx4173, A0=>nx6028, A1=>nx6102);
   ix4188 : or02 port map ( Y=>nx4187, A0=>nx6022, A1=>nx6110);
   ix1859 : mux21 port map ( Y=>nx1858, A0=>LFSROUT_13, A1=>B(13), S0=>
      nx6010);
   ix4210 : or02 port map ( Y=>nx4209, A0=>nx6124, A1=>nx5974);
   ix2101 : mux21 port map ( Y=>nx2100, A0=>LFSROUT_30, A1=>A(14), S0=>
      nx6010);
   ix3837 : nor02ii port map ( Y=>nx3836, A0=>nx6124, A1=>MAC0_MultB_0);
   ix4222 : or02 port map ( Y=>nx4221, A0=>nx6114, A1=>nx6018);
   ix4230 : or02 port map ( Y=>nx4229, A0=>nx6106, A1=>nx6030);
   ix4238 : or02 port map ( Y=>nx4237, A0=>nx6098, A1=>nx6038);
   ix4248 : or02 port map ( Y=>nx4247, A0=>nx6090, A1=>nx6046);
   ix4256 : or02 port map ( Y=>nx4255, A0=>nx6084, A1=>nx6054);
   ix4266 : or02 port map ( Y=>nx4265, A0=>nx6074, A1=>nx6062);
   ix4274 : or02 port map ( Y=>nx4273, A0=>nx6066, A1=>nx6070);
   ix4284 : or02 port map ( Y=>nx4283, A0=>nx6060, A1=>nx6080);
   ix4294 : or02 port map ( Y=>nx4293, A0=>nx6050, A1=>nx6086);
   ix4302 : or02 port map ( Y=>nx4301, A0=>nx6044, A1=>nx6094);
   ix4312 : or02 port map ( Y=>nx4311, A0=>nx6034, A1=>nx6102);
   ix4320 : or02 port map ( Y=>nx4319, A0=>nx6028, A1=>nx6110);
   ix4334 : or02 port map ( Y=>nx4333, A0=>nx6022, A1=>nx6118);
   ix2035 : mux21 port map ( Y=>nx2034, A0=>LFSROUT_14, A1=>B(14), S0=>
      nx6010);
   ix4358 : or02 port map ( Y=>nx4357, A0=>nx6132, A1=>nx5974);
   ix2293 : mux21 port map ( Y=>nx2292, A0=>LFSROUT_31, A1=>A(15), S0=>
      nx6010);
   ix3825 : nor02ii port map ( Y=>nx3824, A0=>nx6132, A1=>MAC0_MultB_0);
   ix4372 : or02 port map ( Y=>nx4371, A0=>nx6124, A1=>nx6018);
   ix4380 : or02 port map ( Y=>nx4379, A0=>nx6114, A1=>nx6032);
   ix4390 : or02 port map ( Y=>nx4389, A0=>nx6106, A1=>nx6040);
   ix4398 : or02 port map ( Y=>nx4397, A0=>nx6098, A1=>nx6048);
   ix4408 : or02 port map ( Y=>nx4407, A0=>nx6090, A1=>nx6056);
   ix4416 : or02 port map ( Y=>nx4415, A0=>nx6084, A1=>nx6062);
   ix4426 : or02 port map ( Y=>nx4425, A0=>nx6076, A1=>nx6070);
   ix4434 : or02 port map ( Y=>nx4433, A0=>nx6066, A1=>nx6080);
   ix4444 : or02 port map ( Y=>nx4443, A0=>nx6060, A1=>nx6086);
   ix4454 : or02 port map ( Y=>nx4453, A0=>nx6052, A1=>nx6094);
   ix4462 : or02 port map ( Y=>nx4461, A0=>nx6044, A1=>nx6102);
   ix4472 : or02 port map ( Y=>nx4471, A0=>nx6036, A1=>nx6110);
   ix4482 : or02 port map ( Y=>nx4481, A0=>nx6028, A1=>nx6120);
   ix4496 : or02 port map ( Y=>nx4495, A0=>nx6022, A1=>nx6128);
   ix2223 : mux21 port map ( Y=>nx2222, A0=>LFSROUT_15, A1=>B(15), S0=>
      nx6010);
   ix4520 : or02 port map ( Y=>nx4519, A0=>nx6132, A1=>nx6018);
   ix4528 : or02 port map ( Y=>nx4527, A0=>nx6124, A1=>nx6032);
   ix4538 : or02 port map ( Y=>nx4537, A0=>nx6114, A1=>nx6040);
   ix4548 : or02 port map ( Y=>nx4547, A0=>nx6106, A1=>nx6048);
   ix4558 : or02 port map ( Y=>nx4557, A0=>nx6098, A1=>nx6056);
   ix4568 : or02 port map ( Y=>nx4567, A0=>nx6090, A1=>nx6062);
   ix4578 : or02 port map ( Y=>nx4577, A0=>nx6084, A1=>nx6070);
   ix4588 : or02 port map ( Y=>nx4587, A0=>nx6076, A1=>nx6080);
   ix4598 : or02 port map ( Y=>nx4597, A0=>nx6068, A1=>nx6086);
   ix4608 : or02 port map ( Y=>nx4607, A0=>nx6060, A1=>nx6094);
   ix4618 : or02 port map ( Y=>nx4617, A0=>nx6052, A1=>nx6102);
   ix4628 : or02 port map ( Y=>nx4627, A0=>nx6044, A1=>nx6110);
   ix4638 : or02 port map ( Y=>nx4637, A0=>nx6036, A1=>nx6120);
   ix4648 : or02 port map ( Y=>nx4647, A0=>nx6028, A1=>nx6128);
   ix4652 : or02 port map ( Y=>nx4651, A0=>nx6022, A1=>nx6136);
   ix4678 : or02 port map ( Y=>nx4677, A0=>nx6132, A1=>nx6032);
   ix4684 : or02 port map ( Y=>nx4683, A0=>nx6124, A1=>nx6040);
   ix4690 : or02 port map ( Y=>nx4689, A0=>nx6114, A1=>nx6048);
   ix4696 : or02 port map ( Y=>nx4695, A0=>nx6108, A1=>nx6056);
   ix4702 : or02 port map ( Y=>nx4701, A0=>nx6098, A1=>nx6064);
   ix4708 : or02 port map ( Y=>nx4707, A0=>nx6092, A1=>nx6072);
   ix4714 : or02 port map ( Y=>nx4713, A0=>nx6084, A1=>nx6080);
   ix4720 : or02 port map ( Y=>nx4719, A0=>nx6076, A1=>nx6086);
   ix4726 : or02 port map ( Y=>nx4725, A0=>nx6068, A1=>nx6094);
   ix4732 : or02 port map ( Y=>nx4731, A0=>nx6060, A1=>nx6102);
   ix4738 : or02 port map ( Y=>nx4737, A0=>nx6052, A1=>nx6110);
   ix4744 : or02 port map ( Y=>nx4743, A0=>nx6044, A1=>nx6120);
   ix4750 : or02 port map ( Y=>nx4749, A0=>nx6036, A1=>nx6128);
   ix4756 : or02 port map ( Y=>nx4755, A0=>nx6028, A1=>nx6136);
   ix4758 : or03 port map ( Y=>nx4757, A0=>nx5986, A1=>nx6024, A2=>nx6136);
   ix5985 : inv01 port map ( Y=>nx5986, A=>nx2412);
   ix4776 : or02 port map ( Y=>nx4775, A0=>nx6132, A1=>nx6040);
   ix4784 : or02 port map ( Y=>nx4783, A0=>nx6124, A1=>nx6048);
   ix4792 : or02 port map ( Y=>nx4791, A0=>nx6116, A1=>nx6056);
   ix4802 : or02 port map ( Y=>nx4801, A0=>nx6108, A1=>nx6064);
   ix4810 : or02 port map ( Y=>nx4809, A0=>nx6098, A1=>nx6072);
   ix4820 : or02 port map ( Y=>nx4819, A0=>nx6092, A1=>nx6080);
   ix4828 : or02 port map ( Y=>nx4827, A0=>nx6084, A1=>nx6086);
   ix4838 : or02 port map ( Y=>nx4837, A0=>nx6076, A1=>nx6094);
   ix4846 : or02 port map ( Y=>nx4845, A0=>nx6068, A1=>nx6104);
   ix4856 : or02 port map ( Y=>nx4855, A0=>nx6060, A1=>nx6112);
   ix4864 : or02 port map ( Y=>nx4863, A0=>nx6052, A1=>nx6120);
   ix4874 : or02 port map ( Y=>nx4873, A0=>nx6044, A1=>nx6128);
   ix4882 : or02 port map ( Y=>nx4881, A0=>nx6036, A1=>nx6136);
   ix4902 : or02 port map ( Y=>nx4901, A0=>nx6132, A1=>nx6048);
   ix4912 : or02 port map ( Y=>nx4911, A0=>nx6124, A1=>nx6056);
   ix4918 : or02 port map ( Y=>nx4917, A0=>nx6116, A1=>nx6064);
   ix4926 : or02 port map ( Y=>nx4925, A0=>nx6108, A1=>nx6072);
   ix4935 : or02 port map ( Y=>nx4934, A0=>nx6098, A1=>nx6080);
   ix4945 : or02 port map ( Y=>nx4944, A0=>nx6092, A1=>nx6088);
   ix4951 : or02 port map ( Y=>nx4950, A0=>nx6084, A1=>nx6094);
   ix4959 : or02 port map ( Y=>nx4958, A0=>nx6076, A1=>nx6104);
   ix4968 : or02 port map ( Y=>nx4967, A0=>nx6068, A1=>nx6112);
   ix4978 : or02 port map ( Y=>nx4977, A0=>nx6060, A1=>nx6120);
   ix4984 : or02 port map ( Y=>nx4983, A0=>nx6052, A1=>nx6128);
   ix4992 : or02 port map ( Y=>nx4991, A0=>nx6044, A1=>nx6136);
   ix5010 : or02 port map ( Y=>nx5009, A0=>nx6134, A1=>nx6056);
   ix5018 : or02 port map ( Y=>nx5017, A0=>nx6124, A1=>nx6064);
   ix5026 : or02 port map ( Y=>nx5025, A0=>nx6116, A1=>nx6072);
   ix5032 : or02 port map ( Y=>nx5031, A0=>nx6108, A1=>nx6080);
   ix5038 : or02 port map ( Y=>nx5037, A0=>nx6100, A1=>nx6088);
   ix5044 : or02 port map ( Y=>nx5043, A0=>nx6092, A1=>nx6094);
   ix5052 : or02 port map ( Y=>nx5051, A0=>nx6084, A1=>nx6104);
   ix5058 : or02 port map ( Y=>nx5057, A0=>nx6076, A1=>nx6112);
   ix5064 : or02 port map ( Y=>nx5063, A0=>nx6068, A1=>nx6120);
   ix5072 : or02 port map ( Y=>nx5071, A0=>nx6060, A1=>nx6130);
   ix5080 : or02 port map ( Y=>nx5079, A0=>nx6052, A1=>nx6138);
   ix5097 : or02 port map ( Y=>nx5096, A0=>nx6134, A1=>nx6064);
   ix5103 : or02 port map ( Y=>nx5102, A0=>nx6124, A1=>nx6072);
   ix5111 : or02 port map ( Y=>nx5110, A0=>nx6116, A1=>nx6080);
   ix5119 : or02 port map ( Y=>nx5118, A0=>nx6108, A1=>nx6088);
   ix5125 : or02 port map ( Y=>nx5124, A0=>nx6100, A1=>nx6096);
   ix5132 : or02 port map ( Y=>nx5131, A0=>nx6092, A1=>nx6104);
   ix5142 : or02 port map ( Y=>nx5141, A0=>nx6084, A1=>nx6112);
   ix5150 : or02 port map ( Y=>nx5149, A0=>nx6076, A1=>nx6120);
   ix5158 : or02 port map ( Y=>nx5157, A0=>nx6068, A1=>nx6130);
   ix5164 : or02 port map ( Y=>nx5163, A0=>nx6060, A1=>nx6138);
   ix5181 : or02 port map ( Y=>nx5180, A0=>nx6134, A1=>nx6072);
   ix5189 : or02 port map ( Y=>nx5188, A0=>nx6124, A1=>nx6080);
   ix5195 : or02 port map ( Y=>nx5194, A0=>nx6116, A1=>nx6088);
   ix5201 : or02 port map ( Y=>nx5200, A0=>nx6108, A1=>nx6096);
   ix5208 : or02 port map ( Y=>nx5207, A0=>nx6100, A1=>nx6104);
   ix5215 : or02 port map ( Y=>nx5214, A0=>nx6092, A1=>nx6112);
   ix5225 : or02 port map ( Y=>nx5224, A0=>nx6084, A1=>nx6120);
   ix5231 : or02 port map ( Y=>nx5230, A0=>nx6076, A1=>nx6130);
   ix5237 : or02 port map ( Y=>nx5236, A0=>nx6068, A1=>nx6138);
   ix5257 : or02 port map ( Y=>nx5256, A0=>nx6134, A1=>nx6080);
   ix5267 : or02 port map ( Y=>nx5266, A0=>nx6124, A1=>nx6088);
   ix5273 : or02 port map ( Y=>nx5272, A0=>nx6116, A1=>nx6096);
   ix5280 : or02 port map ( Y=>nx5279, A0=>nx6108, A1=>nx6104);
   ix5287 : or02 port map ( Y=>nx5286, A0=>nx6100, A1=>nx6112);
   ix5294 : or02 port map ( Y=>nx5293, A0=>nx6092, A1=>nx6120);
   ix5304 : or02 port map ( Y=>nx5303, A0=>nx6084, A1=>nx6130);
   ix5312 : or02 port map ( Y=>nx5311, A0=>nx6076, A1=>nx6138);
   ix5330 : or02 port map ( Y=>nx5329, A0=>nx6134, A1=>nx6088);
   ix5338 : or02 port map ( Y=>nx5337, A0=>nx6124, A1=>nx6096);
   ix5347 : or02 port map ( Y=>nx5346, A0=>nx6116, A1=>nx6104);
   ix5356 : or02 port map ( Y=>nx5355, A0=>nx6108, A1=>nx6112);
   ix5365 : or02 port map ( Y=>nx5364, A0=>nx6100, A1=>nx6120);
   ix5374 : or02 port map ( Y=>nx5373, A0=>nx6092, A1=>nx6130);
   ix5384 : or02 port map ( Y=>nx5383, A0=>nx6084, A1=>nx6138);
   ix5401 : or02 port map ( Y=>nx5400, A0=>nx6134, A1=>nx6096);
   ix5407 : or02 port map ( Y=>nx5406, A0=>nx6124, A1=>nx6104);
   ix5413 : or02 port map ( Y=>nx5412, A0=>nx6116, A1=>nx6112);
   ix5419 : or02 port map ( Y=>nx5418, A0=>nx6108, A1=>nx6120);
   ix5425 : or02 port map ( Y=>nx5424, A0=>nx6100, A1=>nx6130);
   ix5431 : or02 port map ( Y=>nx5430, A0=>nx6092, A1=>nx6138);
   ix5448 : or02 port map ( Y=>nx5447, A0=>nx6134, A1=>nx6104);
   ix5456 : or02 port map ( Y=>nx5455, A0=>nx6124, A1=>nx6112);
   ix5464 : or02 port map ( Y=>nx5463, A0=>nx6116, A1=>nx6120);
   ix5472 : or02 port map ( Y=>nx5471, A0=>nx6108, A1=>nx6130);
   ix5478 : or02 port map ( Y=>nx5477, A0=>nx6100, A1=>nx6138);
   ix5498 : or02 port map ( Y=>nx5497, A0=>nx6134, A1=>nx6112);
   ix5508 : or02 port map ( Y=>nx5507, A0=>nx6124, A1=>nx6120);
   ix5514 : or02 port map ( Y=>nx5513, A0=>nx6116, A1=>nx6130);
   ix5522 : or02 port map ( Y=>nx5521, A0=>nx6108, A1=>nx6138);
   ix5540 : or02 port map ( Y=>nx5539, A0=>nx6134, A1=>nx6120);
   ix5548 : or02 port map ( Y=>nx5547, A0=>nx6126, A1=>nx6130);
   ix5556 : or02 port map ( Y=>nx5555, A0=>nx6116, A1=>nx6138);
   ix5573 : or02 port map ( Y=>nx5572, A0=>nx6134, A1=>nx6130);
   ix5579 : or02 port map ( Y=>nx5578, A0=>nx6126, A1=>nx6138);
   ix2310 : mux21 port map ( Y=>nx2309, A0=>nx4766, A1=>MISR_out_30, S0=>
      nx6010);
   ix4767 : xor2 port map ( Y=>nx4766, A0=>RegOut_dup0_30, A1=>MISR_out_31);
   ix5606 : or02 port map ( Y=>nx5605, A0=>nx6134, A1=>nx6138);
   ix2300 : mux21 port map ( Y=>nx2299, A0=>nx4760, A1=>MISR_out_31, S0=>
      nx6010);
   ix4761 : xor2 port map ( Y=>nx4760, A0=>RegOut_dup0_31, A1=>MISR_out_0);
   ix4567 : oai32 port map ( Y=>nx4566, A0=>nx6134, A1=>nx6138, A2=>nx5988, 
      B0=>nx5602, B1=>nx5990);
   ix5987 : inv01 port map ( Y=>nx5988, A=>nx4536);
   ix5989 : inv01 port map ( Y=>nx5990, A=>nx4538);
   ix2290 : mux21 port map ( Y=>nx2289, A0=>nx4754, A1=>MISR_out_0, S0=>
      nx6010);
   ix4755 : xor2 port map ( Y=>nx4754, A0=>RegOut_dup0_0, A1=>MISR_out_1);
   ix2280 : mux21 port map ( Y=>nx2279, A0=>nx4748, A1=>MISR_out_1, S0=>
      nx6010);
   ix4749 : xor2 port map ( Y=>nx4748, A0=>RegOut_dup0_1, A1=>MISR_out_2);
   ix2270 : mux21 port map ( Y=>nx2269, A0=>nx4742, A1=>MISR_out_2, S0=>
      nx6010);
   ix4743 : xor2 port map ( Y=>nx4742, A0=>RegOut_dup0_2, A1=>MISR_out_3);
   ix2260 : mux21 port map ( Y=>nx2259, A0=>nx4736, A1=>MISR_out_3, S0=>
      nx6010);
   ix4737 : xor2 port map ( Y=>nx4736, A0=>RegOut_dup0_3, A1=>MISR_out_4);
   ix2250 : mux21 port map ( Y=>nx2249, A0=>nx4730, A1=>MISR_out_4, S0=>
      nx6010);
   ix4731 : xor2 port map ( Y=>nx4730, A0=>RegOut_dup0_4, A1=>MISR_out_5);
   ix2240 : mux21 port map ( Y=>nx2239, A0=>nx4724, A1=>MISR_out_5, S0=>
      nx6012);
   ix4725 : xor2 port map ( Y=>nx4724, A0=>RegOut_dup0_5, A1=>MISR_out_6);
   ix2230 : mux21 port map ( Y=>nx2229, A0=>nx4718, A1=>MISR_out_6, S0=>
      nx6012);
   ix4719 : xor2 port map ( Y=>nx4718, A0=>RegOut_dup0_6, A1=>MISR_out_7);
   ix2220 : mux21 port map ( Y=>nx2219, A0=>nx4712, A1=>MISR_out_7, S0=>
      nx6012);
   ix4713 : xor2 port map ( Y=>nx4712, A0=>RegOut_dup0_7, A1=>MISR_out_8);
   ix2210 : mux21 port map ( Y=>nx2209, A0=>nx4706, A1=>MISR_out_8, S0=>
      nx6012);
   ix4707 : xor2 port map ( Y=>nx4706, A0=>RegOut_dup0_8, A1=>MISR_out_9);
   ix2200 : mux21 port map ( Y=>nx2199, A0=>nx4700, A1=>MISR_out_9, S0=>
      nx6012);
   ix4701 : xor2 port map ( Y=>nx4700, A0=>RegOut_dup0_9, A1=>MISR_out_10);
   ix2190 : mux21 port map ( Y=>nx2189, A0=>nx4694, A1=>MISR_out_10, S0=>
      nx6012);
   ix4695 : xor2 port map ( Y=>nx4694, A0=>RegOut_dup0_10, A1=>MISR_out_11);
   ix2180 : mux21 port map ( Y=>nx2179, A0=>nx4688, A1=>MISR_out_11, S0=>
      nx6012);
   ix4689 : xor2 port map ( Y=>nx4688, A0=>RegOut_dup0_11, A1=>MISR_out_12);
   ix2170 : mux21 port map ( Y=>nx2169, A0=>nx4682, A1=>MISR_out_12, S0=>
      nx6012);
   ix4683 : xor2 port map ( Y=>nx4682, A0=>RegOut_dup0_12, A1=>MISR_out_13);
   ix2160 : mux21 port map ( Y=>nx2159, A0=>nx4676, A1=>MISR_out_13, S0=>
      nx6012);
   ix4677 : xor2 port map ( Y=>nx4676, A0=>RegOut_dup0_13, A1=>MISR_out_14);
   ix2150 : mux21 port map ( Y=>nx2149, A0=>nx4670, A1=>MISR_out_14, S0=>
      nx6012);
   ix4671 : xor2 port map ( Y=>nx4670, A0=>RegOut_dup0_14, A1=>MISR_out_15);
   ix2140 : mux21 port map ( Y=>nx2139, A0=>nx4664, A1=>MISR_out_15, S0=>
      nx6012);
   ix4665 : xor2 port map ( Y=>nx4664, A0=>RegOut_dup0_15, A1=>MISR_out_16);
   ix2130 : mux21 port map ( Y=>nx2129, A0=>nx4658, A1=>MISR_out_16, S0=>
      nx6012);
   ix4659 : xor2 port map ( Y=>nx4658, A0=>RegOut_dup0_16, A1=>MISR_out_17);
   ix2120 : mux21 port map ( Y=>nx2119, A0=>nx4652, A1=>MISR_out_17, S0=>
      nx6012);
   ix4653 : xor2 port map ( Y=>nx4652, A0=>RegOut_dup0_17, A1=>MISR_out_18);
   ix2110 : mux21 port map ( Y=>nx2109, A0=>nx4646, A1=>MISR_out_18, S0=>
      nx6012);
   ix4647 : xor2 port map ( Y=>nx4646, A0=>RegOut_dup0_18, A1=>MISR_out_19);
   ix2100 : mux21 port map ( Y=>nx2099, A0=>nx4640, A1=>MISR_out_19, S0=>
      nx6012);
   ix4641 : xor2 port map ( Y=>nx4640, A0=>nx5633, A1=>nx5733);
   ix5734 : xor2 port map ( Y=>nx5733, A0=>RegOut_dup0_19, A1=>nx5782);
   ix2090 : mux21 port map ( Y=>nx2089, A0=>nx4632, A1=>MISR_out_20, S0=>
      nx6014);
   ix4633 : xor2 port map ( Y=>nx4632, A0=>RegOut_dup0_20, A1=>MISR_out_21);
   ix2080 : mux21 port map ( Y=>nx2079, A0=>nx4626, A1=>MISR_out_21, S0=>
      nx6014);
   ix4627 : xor2 port map ( Y=>nx4626, A0=>RegOut_dup0_21, A1=>MISR_out_22);
   ix2070 : mux21 port map ( Y=>nx2069, A0=>nx4620, A1=>MISR_out_22, S0=>
      nx6014);
   ix4621 : xor2 port map ( Y=>nx4620, A0=>RegOut_dup0_22, A1=>MISR_out_23);
   ix2060 : mux21 port map ( Y=>nx2059, A0=>nx4614, A1=>MISR_out_23, S0=>
      nx6014);
   ix4615 : xor2 port map ( Y=>nx4614, A0=>RegOut_dup0_23, A1=>MISR_out_24);
   ix2050 : mux21 port map ( Y=>nx2049, A0=>nx4608, A1=>MISR_out_24, S0=>
      nx6014);
   ix4609 : xor2 port map ( Y=>nx4608, A0=>nx5633, A1=>nx5758);
   ix2040 : mux21 port map ( Y=>nx2039, A0=>nx4600, A1=>MISR_out_25, S0=>
      nx6014);
   ix4601 : xor2 port map ( Y=>nx4600, A0=>nx5633, A1=>nx5763);
   ix5764 : xor2 port map ( Y=>nx5763, A0=>RegOut_dup0_25, A1=>nx5780);
   ix2030 : mux21 port map ( Y=>nx2029, A0=>nx4592, A1=>MISR_out_26, S0=>
      nx6014);
   ix4593 : xor2 port map ( Y=>nx4592, A0=>RegOut_dup0_26, A1=>MISR_out_27);
   ix2020 : mux21 port map ( Y=>nx2019, A0=>nx4586, A1=>MISR_out_27, S0=>
      nx6014);
   ix4587 : xor2 port map ( Y=>nx4586, A0=>RegOut_dup0_27, A1=>MISR_out_28);
   ix2010 : mux21 port map ( Y=>nx2009, A0=>nx4580, A1=>MISR_out_28, S0=>
      nx6014);
   ix4581 : xor2 port map ( Y=>nx4580, A0=>RegOut_dup0_28, A1=>MISR_out_29);
   ix4801 : and04 port map ( Y=>nx4800, A0=>MISR_out_26, A1=>nx5992, A2=>
      nx5753, A3=>MISR_out_23);
   ix5991 : inv01 port map ( Y=>nx5992, A=>MISR_out_25);
   ix5785 : nand04 port map ( Y=>nx5784, A0=>nx5743, A1=>nx5738, A2=>
      MISR_out_20, A3=>nx5728);
   ix5787 : or04 port map ( Y=>nx5786, A0=>nx5723, A1=>nx5718, A2=>nx5713, 
      A3=>nx5708);
   ix4839 : and04 port map ( Y=>nx4838, A0=>nx5703, A1=>nx5698, A2=>nx5693, 
      A3=>nx5688);
   ix4849 : and04 port map ( Y=>nx4848, A0=>nx5683, A1=>nx5678, A2=>
      MISR_out_8, A3=>MISR_out_7);
   ix4861 : and04 port map ( Y=>nx4860, A0=>MISR_out_6, A1=>MISR_out_5, A2=>
      nx5653, A3=>nx5648);
   ix4871 : nor04 port map ( Y=>nx4870, A0=>nx5643, A1=>nx5638, A2=>
      MISR_out_0, A3=>nx5994);
   ix5993 : inv01 port map ( Y=>nx5994, A=>nx2335);
   ix5995 : inv01 port map ( Y=>nx5996, A=>nx2347);
   ix5997 : inv02 port map ( Y=>nx5998, A=>nx5996);
   ix5999 : inv02 port map ( Y=>nx6000, A=>nx5996);
   ix6001 : inv02 port map ( Y=>nx6002, A=>nx5996);
   ix6003 : inv02 port map ( Y=>nx6004, A=>nx5996);
   ix6005 : inv02 port map ( Y=>nx6006, A=>nx5996);
   ix6007 : inv02 port map ( Y=>nx6008, A=>nx5996);
   ix6009 : inv02 port map ( Y=>nx6010, A=>nx5996);
   ix6011 : inv02 port map ( Y=>nx6012, A=>nx5996);
   ix6013 : inv02 port map ( Y=>nx6014, A=>nx5996);
   ix6015 : inv01 port map ( Y=>nx6016, A=>nx5848);
   ix6017 : inv01 port map ( Y=>nx6018, A=>nx5848);
   ix6019 : inv02 port map ( Y=>nx6020, A=>nx5844);
   ix6021 : inv02 port map ( Y=>nx6022, A=>nx5844);
   ix6023 : inv02 port map ( Y=>nx6024, A=>nx5844);
   ix6025 : inv01 port map ( Y=>nx6026, A=>nx5864);
   ix6027 : inv01 port map ( Y=>nx6028, A=>nx5864);
   ix6029 : inv01 port map ( Y=>nx6030, A=>nx5860);
   ix6031 : inv01 port map ( Y=>nx6032, A=>nx5860);
   ix6033 : inv01 port map ( Y=>nx6034, A=>nx5872);
   ix6035 : inv01 port map ( Y=>nx6036, A=>nx5872);
   ix6037 : inv01 port map ( Y=>nx6038, A=>nx5868);
   ix6039 : inv01 port map ( Y=>nx6040, A=>nx5868);
   ix6041 : inv01 port map ( Y=>nx6042, A=>nx5880);
   ix6043 : inv01 port map ( Y=>nx6044, A=>nx5880);
   ix6045 : inv01 port map ( Y=>nx6046, A=>nx5876);
   ix6047 : inv01 port map ( Y=>nx6048, A=>nx5876);
   ix6049 : inv01 port map ( Y=>nx6050, A=>nx5888);
   ix6051 : inv01 port map ( Y=>nx6052, A=>nx5888);
   ix6053 : inv01 port map ( Y=>nx6054, A=>nx5884);
   ix6055 : inv01 port map ( Y=>nx6056, A=>nx5884);
   ix6057 : inv01 port map ( Y=>nx6058, A=>nx5896);
   ix6059 : inv01 port map ( Y=>nx6060, A=>nx5896);
   ix6061 : inv01 port map ( Y=>nx6062, A=>nx5892);
   ix6063 : inv01 port map ( Y=>nx6064, A=>nx5892);
   ix6065 : inv01 port map ( Y=>nx6066, A=>nx5904);
   ix6067 : inv01 port map ( Y=>nx6068, A=>nx5904);
   ix6069 : inv01 port map ( Y=>nx6070, A=>nx5900);
   ix6071 : inv01 port map ( Y=>nx6072, A=>nx5900);
   ix6073 : inv01 port map ( Y=>nx6074, A=>nx5912);
   ix6075 : inv01 port map ( Y=>nx6076, A=>nx5912);
   ix6077 : inv01 port map ( Y=>nx6078, A=>nx5908);
   ix6079 : inv01 port map ( Y=>nx6080, A=>nx5908);
   ix6081 : inv01 port map ( Y=>nx6082, A=>nx5920);
   ix6083 : inv01 port map ( Y=>nx6084, A=>nx5920);
   ix6085 : inv01 port map ( Y=>nx6086, A=>nx5916);
   ix6087 : inv01 port map ( Y=>nx6088, A=>nx5916);
   ix6089 : inv01 port map ( Y=>nx6090, A=>nx5928);
   ix6091 : inv01 port map ( Y=>nx6092, A=>nx5928);
   ix6093 : inv01 port map ( Y=>nx6094, A=>nx5924);
   ix6095 : inv01 port map ( Y=>nx6096, A=>nx5924);
   ix6097 : inv01 port map ( Y=>nx6098, A=>nx5936);
   ix6099 : inv01 port map ( Y=>nx6100, A=>nx5936);
   ix6101 : inv01 port map ( Y=>nx6102, A=>nx5932);
   ix6103 : inv01 port map ( Y=>nx6104, A=>nx5932);
   ix6105 : inv01 port map ( Y=>nx6106, A=>nx5944);
   ix6107 : inv01 port map ( Y=>nx6108, A=>nx5944);
   ix6109 : inv01 port map ( Y=>nx6110, A=>nx5940);
   ix6111 : inv01 port map ( Y=>nx6112, A=>nx5940);
   ix6113 : inv01 port map ( Y=>nx6114, A=>nx5952);
   ix6115 : inv01 port map ( Y=>nx6116, A=>nx5952);
   ix6117 : inv01 port map ( Y=>nx6118, A=>nx5948);
   ix6119 : inv01 port map ( Y=>nx6120, A=>nx5948);
   ix6121 : inv01 port map ( Y=>nx6122, A=>nx5960);
   ix6123 : inv01 port map ( Y=>nx6124, A=>nx5960);
   ix6125 : inv01 port map ( Y=>nx6126, A=>nx5960);
   ix6127 : inv01 port map ( Y=>nx6128, A=>nx5956);
   ix6129 : inv01 port map ( Y=>nx6130, A=>nx5956);
   ix6131 : inv01 port map ( Y=>nx6132, A=>nx5968);
   ix6133 : inv01 port map ( Y=>nx6134, A=>nx5968);
   ix6135 : inv01 port map ( Y=>nx6136, A=>nx5964);
   ix6137 : inv01 port map ( Y=>nx6138, A=>nx5964);
   ix6139 : inv02 port map ( Y=>nx6140, A=>MAC0_MultB_0);
end Behavioral ;

